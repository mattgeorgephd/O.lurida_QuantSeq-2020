�      ��[�&�q�	��6q$H����)P�D���RU�KU��Y};k����Ew�8�A�UO�'_���턔��SΈp��k���������~����fU�X/��B���?��/�������z��~�������_�����������������?�?U/�_/|����O���������'�ۿ�����^�l�S���X�޵������k�U����������.m���w�qi���M�[m���������m��ʓ~��wv��-Ow�K��j�z�<�q�����߿t~�6����|wi{��_[|<�x��wi�z|�����o���a��jy.oM�kۃϻ��w�|������=�j�����|��˥����sm>|h���w绶~�������?4<t�?o�k�s����7�ί��?�[=���q�>6?���_Z�km�X?g�w�z��u�_��j�ϖ��ϛ�V����翶���.Ϳg���Ʃ�|���C��|���E�l�������������k���ޗ��k�˥�wi~=��i�|��������<�^���������}��9{������|M�k�[��K����?t����6����w]�_����yW�k�~ߴ�������ۇ6��&����_��_Z>[��m���?{��并��}\�������_�߯��CS�o�����������b띭?߷��Z�k�{��ϛ>g�m<~��I��o����|��GW���|���Z��������ǵ���l|m�_z��͟׎�t����cӇϿ����o�|���g�wv<?4�W�����v���][�oZ�;{�K�ߥ�Y-_w����|}���ϟ7|��ߗ������m��4������g�=��l|�=V�w�x���]y��޵�͵ǩ�����X����^:]Z�k�S}���~���������7����^��c����c�򟭿Ϳz�K�mW���?��������f���?��_�������^*������ז�y�����/�������jy9_w�k�w���������C��y����^�����>�OΖ���s�}�^?���|�Z���O�����{����m�<4~�6�>�qW_>���o����?4�|�Ǵ��Wۿ�޵�����C���&�9[�k�������>��si{\�O�����]}�|�׿v<����[-�C�~����}ܵϥ�����w�{�����]{|i�l����=�|v6޺�_�>6�j���?{���?��s6_]�����_��Ζ���z��硭����_:�4�]�_�}�����C�׫�_�߇n�T���=��j}�������>���k˷�_����ׇn�k�g�u�K��ʳ�>��o��g?�����]��{>��z����Cϗ���;_�����m��.�j�������i�a�|��g�w�|���}���<�������q��}L�M���k�w�x��<g�;?t~}���s_��׶���ؕ�y���>6���/�������>4�<���w?�c��=?�?��}����������ז����ٟ�W�wm�_-���l{t�?;�?��.=�}�����K�����-�7m����|6^���.�wg�۝/������_[���O��q�m�k���w�z������������C�����l���]�Z�?�|�Z߮=��8{������l<������|�����qW����_W�t���=[�K���忶���׶��󟍿K�����=N�M���?�|u��q�|�?o�����t|m����_;_������'������񸚟~^��K���_=���w绶?.��K�9����j�W�k�oߧ�w�[���揳�٥�s�����y_[�t���6�t>�t�^m��|�]���66�p|m�.����?4{\/��y��^<����qw���<��j}������}h�k�g�w�����{h�=o����g��������۝Ͼ_-��]&ϥ�����H�[�~�������M�{m���/-/�{h�v���������t�?[��ϛ<��o����']���^;�/=6�R����7{_�M��}���߳����o��=~ژ�u��ηz�K����}�Z���s�[��������?�_�^:�����g�������=��&o:W�������ٗ������w��g����O���l�����{���=�7M޳�_=w>~�|����]?��O�;������������ɿZ�K��}�;�j�����ߵ���?4�/��7M�k���M�K��տ����t��������][��6���}����=l|m}ژ���������K�-��_;~��M���={��>~h���-���9��ߵ�����>��,��^�l{��_[_�o㇦O*��6~�|��]y��w�>Mއ���m�M��y��K�������=�c�z��������<M�t���?�{?������=���ўw����������]5�.=���m|m{=�q�߷���]�~������v|>�������;���^[��}���߫׻���^�락���;[_��l}M�k�����ك���������֧+�_Z�K�%��l{\Z�k�{m�^z�k��C����\{��M�����6ߵ�=�~�������l�/=��j�l��|�彴=�����u�{h�_:V�;�����׻t���m|m�\;^�=���y�~g�����]�y�������o�~���j�����N�=[����|g�z�K�����g����{h���w��M����oڸ����z�^�l�S���8��k����I�h��C���Ζ���=�?��{�㮾������]�߫�;��彶�.-��66��W�m�����W����m�n<��OW���<o���s���?���-�C�����ƴ�m�����.�����|~�}V�ߕ���Y-��~�=Ζ��f�k��|��]y����z��϶o�>����_�]����k�M�T��f����|����ϖ��_���}��z2�}��9�7yL�t>�����M�����S��}Wo������7��=O����=���U�3�|\�㮾����_�O���3}����/�����_��x���O��ߧ����x��+壳����yu>��Q����]�(_��ή�R~;���x[�-���g:���x��S�����M��T���I:�zw�������է�'������٥�_���|��su}�շ�Ƿ]<��W����F{v���u�:R}��]���0�t�ڍ��>�t>������^ZO����]�R���ש<i��x������x���)~R{����_��g���꟮ߕ?�G7�����˪^�x�����|�W������j������]�����o]~�ړ�v����ɓ�#��������t�Ѝ���:��j~����z���jw�������������ǵ�|&��m���Wק��"�g�_��]����xK���}6?��7l�n�ٍ��~}��]{u�Ϫ��aϻ�t�۵��������?�������|���墳(o������u�c��C�WU���F�Vۯ�o�z��L�?�|u���������������_�|�Ow?��7�k���|��Kj�ԟ]�t����i���oi}�Z����]~��-��4����k:N�]����׍�n=h�3{�z�~u����]��c�'�w7���N�~ߵg7^ζ7�S�����������K�'�����|׎������j��g���y7>;�qO��oi�>۟�������jUVo�y��V??��~6^��H�K�_]�>W�gR���GV���z������������_*�O��Ϳ]�w�{6��u�׍���0]�������k���K���������e���������J������7��*�G�x?�J�/�i�v���׎�?��C7^h��>������s��I���>;�]��������g�����_�����^\]?�ݟ9����G��*�[����1�]��\�W��V�i5\;����UY���S����i������[�?�x�=9��qu~N��Ξ�˯6:>{���o���g�)��O���M���|��ʻ����V����?���w�M����t�7������������_V�'���7�w�||��_>�zbu���_����#���?_]~��OW����ڞ\�޷��x�Η�?�g_�}�����u*��x6�]��:�R��>g��j�R~�S�����4���j�V������2y������u�)�K�W燔?��|U��W�W���|}�>�����ou��Ń��������^���n�����~��z�]}(_�?�����|wv|����1]�[_�����(��S�V��]�u���߮�R{r�����sw�Ծi�������Q��֧g��L�n~����]?]}��M������z��T����ڷ��K���[UV�v�����p�7\ou<w���?�G����R��K˟����WV���êl?�Z�/]���7�/�7���Տcʛ�W��L�K�]�2y���|g믮���_z?q6~�z��j�������[_��w���z4��k���e�VϷz�B{���n�p6_����|ѝ�*���������J���w6_t���EU���������>����şɛ�������j�������Cw���j���T���L�w6���oо�����&���ߍ��|��Ծi��]?Ue��������z���H�7�����Iw��Z��_�x��3��<��xN���ou��և]�t����3շ������^i���g�V��]}����]W�Կ�z��R>8{���3���o�O�����z��g������Ryh�������5���l�t���~Z?���~W�n���Q�ۯ�x��3�O��Jמ���v�}vc5^���j�t��ѵg�]���3����'���>|�|���]�����;�j~[]?Ӟf߮|����˴��|������~]|��k�_��Y]?��<�~)���.~��X-���u����ݏu��gg���z�l����C�O�g��_����6>_�����]<t�!�g�~]<t���g�����﫲�u�yj�׭/�x8��@}W�׵g7�v���8�o*�ً�w���ߝ���/�?��˟�z����w���w6�T����|�[^��խ��󙼴o��k?��[߭��l����������~U�{����Z�oH�K���}����k��W��t�ѵO:j�tӵ��)����jcʗ���ǥ�|u}ۍ��,?t���'ζ���ԟi<We���c����K����N���;�?��]{����xh����qW�T_���C�^����'�o5?��&�7�^�~)����j>Z�?��g�=�ϥ�ǫ�+O:w��������|l�w�pu~7����u�����)���G�_��ד��Y�����}oc���Mӏߧ��x�}����o���ll�v��ʗ�:ޫz��ƫ�)_�O[5��,��xN�8կk?��凳񑎻���G�]<t��sW?�v=ҵw7\{�._w���wU����[?������g׋�^�oή/L�Ԟ]��]?��g��_��ҭ�(o�_i�r��"�?�u�zju����Rj�ʏg�'էˇ]{���������~�?�|a������G��g�ˇg�o���������8����ϳ��]{v�����U���u�Wg�;��j����|i�W�w�}��ӭWϷ�~�zn����z���gu>>ϫ����ѭ��x<;�W��4�xN�E�W�ow�~o�X���z�������[��񼺿v6���_^]t��[��������ɳ_U߮��t���wu}٭��}>_ϫ����n��t�]u��n�>������[u�_m_�[u�g�C���.�S�����+�z��_���>﮿�UY`5�\{tm���?��}��������ҝ?��W�����\�l~���K�[����M���㹻��[���n�nc�߮�������.��������7f>_]Ϭ�ov���x�������^�x1{��O�zc���뛽R�����=��J7��&�W����x]m��>]���=;�V�'��L�._w�n㴞�t��z����|���^�jm�v뿳������_]O��S����l�u�c�i~��W�?�����S����j���n�����||��V׷�~�l���7S�4}-?t�[�_]m����������y��j}W��j|�ο��Pu������Ky��٭_Wۯ[ow�{��OW㽛V�W����t>M�������������ݟ����9�������Nj��l���ӭ�.͗���������n|��O��&�Og���O�:��o�}Z�<�K�;������+�zau���6��������_]o�]?��W��Ϭ��ls�����pj�n���I����������ЭO�����~Z/v�(���ϻ��n>�֧���K�׭W/�0~����~"�3�4�R��Fw?ѭV�OL�����t��Z����;��<�g��i=qv=حV˓��^��#]|�������x]]�X}v6��������]}W˟���|��Gu�$�7�������ܕg5������wv���������IW�����i���ͥ����|���]�ϴ�M�s��ڭw���v�ѭ�������/�׭R{��õ�өV���x���j{��t�{����|�Z�K�Ci}��J��������������z�z��k��]>����#f�4^Ϯ���au�����⽋�������Ⱬ��z�������K�w����������n�Nyή�m}�O��������t?׍?���zi�~2�ww��_�|z�x��3������������ݟ���t������w�W�������گ�O��7ԧk�n����t�n<u�������z?��>����G{r|��ڍ�����֛f�����������ם/������Y����i����_z�vv��������N��t=zv�i�<�~7�x5>(���9���8�'�ۿt~�����������_��?^	����M�3{��8�7�M~ӗ��|�7�'�g���;�W�6?�O�c�|�ڷ�������c�H�9�'�1�R��8�{ʏ�_���.��x4Tm���4ߦc�?�7����m5_����S��c��&j��T���K�S�7>R|ql�^��n�dx��w�|i<�u��|?����~ ��n�ԭ�����u�/�7���w�+��t���C�i����=O��/�����6{��f��������+���Э��|�}?�w�1���g���>�S�X������E�������_���t�!�_�q���w�o���O�]���o�����폤�Nj/�?��n�ݵg���w)���ZW�4���q����]��|i�ۿ���?�z(�5�w�������;���S>L��)����H��?�_*_Z���u���?N㯋����ƿ���M~�/����擴^��M���T�.�t����t��Ҟ����~jZ���`�/�W�|��L�0��4V����.�R�n�w�M���z�{�d�J��#��t�+��������W��j��Y�T�4���n������^N�%��~M�מWe�O����ή��߯Οi�����拴_����|��|n������q�����z���e���U�x��n=b�4>H���S�����t���~���X�~�ֳ��7UY�-���~f����U�N���_V�k����8��ͯf�4~���)�ߺ���p����[���������ٞ��i}��c�/R���J�ww�:^S��~��._t����|޵?�ݭg�����)?��z��?��ϴ����t���'������K�'�O�]�O������~����/��K����s��?]�X|�x�ڷ*����n?=�������_ӷ[?��^�����]����J����=����,>8_��N��i�����ɟ�/է[_�����)?W�������axN�i�u����$�/�'�;��8����ԭ��^J�]�tϧRy����o����m���Q��6>��S~��_�~��SyVׯi=�:�,��oh�4�������ش^L����^��2����n�����Mi�W��'t��i>�ڣ˗�~��~k�U����OH�����[�����[S��)�w�k���|i���C�7ʛڣ�i��:�c�o�n?&����.߬�w�z&�O���������+�����S<u�ii ���t�7�_���<��?�O뇳��ƫɓ����g�\��K�m&��g��I7�������������O��k�����%�_��OUV����?��S~Z]u�u�^�O�]�����i>L�s�������c)�->����/�O7_������q�?Z]��<�~����j���_]���x4<��N��ߍ�t=�w��n��z��}UY}���_w?g�J��[�[=�����!շ˿)^�z�[���ϵ���=S~J�}_|��o�q=���V�{]���Ӵ�����_��4?t���l�n`��g׿����ߴ���o��J�i$��|��ӭ����f���j����� ��n>;��0�Ӟg��t�d�խ���T���i<���ݏ�����|�ͯ]����S�u��i|��[o��U��W�^���yY��t�����/��,�ۭW�|����x2{��7���n>��K]������)�S�J�C����8ŋ�W�~_��Zw?�:����>��gf�n�L�/�����O퓎S�W�S~����M��������I�K���3�O����t?ҍ/�.���&�g��I��{*Oʯ�� ��n���_��)�����x�����m���[�_i��.^S���ܾO��G�tϯ8���)�����H7?�����i~��.~�xM���?���.W�?���ǔ?���|��R>��i?�{`�\��t���]�g��n?��k�u�ۺ��n?�[��t?L�w��i���w����]�-~S~��?R�������L�_�?[mϔ/�x��9^�_i}��������k��I�.��xN�C�g�1�S}��k�H������L�Wڟ3|t�*�o�_�|5?v�;��������Ru\���|؍ߔ_�������:ޭ�4~�������[w�ؕ�긿��Ǥ�Y���?;�X�L�M�i��� �u��������qZϙ}���>f��<f��I�����i}�=X]o������<����K�/i?��?��ߑ��k�K���W�'�}:�����4{�_��^x�<�'�#^_��z�~��S�W��|ߘ�����M���t��7�����6�����g�3��|�[?)�S<������g����;�٫j˷f�?��L~�����i���3��O�)�S>��������c�����4��2}V�']����[u�ֿ�)�u�)�g�Wi�n|��[u�ҭW�����:�oZ��]}R|���?���z7�g�w���:_�������n����������)>�2|��?V��y7����z?����oi"�'g����e�O�|�:~���?����?���~w��ҭ��������'����7~��Q׾]~��ԧj�w����%ū�#�g������c��qW�K���w��S>��#�|d������֭���������/�����F��m=~o�n=�����ϻ����V���:�C�ǫ�x5��->��Hy�����yL*��������S~o�x5���{�~��OH��o�Ϻ��=��é_�����������/W�_���=���N����֫)�|��Kw��ݟt����j}�������j>]�?I��n�����D����|ju����i��^]����������C��~Z�?5��)���z��f|`��M����|��?�|i|mx��n?pu~����S�Z�t�K)�t�s��_מ]~<{����{~q��W��U���4����=OY}���T~���n����z?]?���zuu|v��q������b�J�9��.>��e�Q^��?L�g���?��n�K�O������Mڿ�x���n~_����|7��������?��S>Y�߹^���i������ڧ{���t��?[������?��_��_��0{��#��.����ԟ&��{���'�o��GR>]/�����������Ծ]�����x��K�Q���~�������V�S���˩<�T���>J�)ߛ=��<�?���[���_T�%��ū���_s��?i'����^����������QW��R���_W�n���U�O��ڥ��������H�4�|�z�K����zi�ԭ�R���������γ�K������z8����*�O�������Ot�=���u�5��h��i����|d���$��[O��?��oZ_t�!��b�U����z��~n7�v뛳����ⷻ_M�s6�������?�᩻���F�_���C�����)_�<��w��\��W����n=��n����TޔS���L�O�j�m|�����+�T�.?�����/)�[�ظ�_M���Ol�������oʧ���~=����|����c�[��R>N�;�|�z�j���q�Wi���m�^uO��������]�g����*�G�?�z��1����Ϯ�V�oR�Y�v����j�/���H�?��s*���~O��|c���������[ϧ��3}���T�4�������������$����`5�-��s�?���~0�Z����~i>���,�|ԗ��3Η���~t�~Z?���7�_��[���������9}��%������Ͼ���kw���7��t���ֳ�8�?��̞i}��R�����>���_�/c��z0~�)�x��5���S�}��}���m�;�U^>���9��s�G���|n�0��=߯'k����5{�����gx�|���e��8�3�k����k��s�G���5}l������ƣ�#�3���յǖo8N���_�|a�I���`�N�Q����_�-o�/)��i<�x7>���û�#�O�~K��fÓ�c|��eZ/��_�_�g�_u\ߤ���%�C��4^��i������]���+�����f?���O���h�`��ˇi�u��t?��{����֋�~��w�a�k�[�'�O��O��\��4���@ʧ�_�q~N�w������������z���%�/�/�gi=������y����{��AZ��=R�7>I�)�����n�I��W���c>N�/)���lx��i���_J����*���D�O��H���q��T���Jڏ㸻J�#��@�~�O�����W��6~I�ۏ���t}��Oi}����Kzސ��~T�~���O��}���[|?���m|�����i�,ݯ��<�n?��gi��փ)����~>w�;��=O�ֻ&O�^�<��a�����g�O��7���˴�J���w��t���������R~L��,?u���Q���)^�����m�o�?�z�ۯ2���xI�[V/����^�� �M�C������͟�~(�*_/�'��x�ֳ)���o��'=����������W�o�O�o�����׭__�|]<��۴>%^�{?�[˧i�Fy�xJ�O�;��4���C���������m������������]��A�i?:�7�����H�O������"�O�G�GV���8�W�OY����:������sz�#�o�=��_���?�Ǥ���&�����?�ߥ�|��CZ��yH��M�a��5<�}��K�[_�~���<ݏ��z�?O�Sʛ�R�H���o��i>����־O�I����}�+���������.���핮��O�|���Dw���oX|��T�O���1�ϲ���'���������ɳ�o���/=?O����/=/��=��~N�?ګ{�'�[�7˟�y��n�I�mi�tσR�����W��i��[��?��J�o�Ou�����w��/�?V������3h���S�Y?9埴~螇���4����t�֭��<�/��f�'���|_����O����|����"���M���~:=��z'}�+_��1퇦�tʿ�}�|,��S>�:��n�=�_�_��Ξ�w�i����n?(���S���Kw������Dz���cR|�����l�w�M����#폙���3�/��ƣ�_u|~d������-���o����&����u뿴�1�̿)t�O-����켺���}j�K�Kw��=I���O��� �w��i=c�K��cߧ����6�L޴��|�?�������>M�+�Wm?i|��_���Կi<t���?i>H�����<��s�����n���S����S{���/�8���Ϧ������~��7��Z|���i~K�Ai=���{^L{�����?��Ԟi���of���Z�ǜݿH���(��i�I�M�W�������~j�?R��<��_�y��Կ��V���M�gS��xK���_�o7������f��yL�<�g�/�z3���U�����c/��{���4�����_�~��c��n��:ߥ�����4w׻t�f��[����*돧����n���1����I*O�_�=?랯u��n��[?Z>H�7��g�o��k��zz�=��}���o����a�����W��Y]�����/��|����_��X��8�g�_��L�5[��8��u�櫪��䴾L�gگN�c��4���R>N���<�s���]�G6�?��x��b�M�#�ʟƋ���=��?D3������������j��_:���o���>�\�����=�^=yg���?���o�������ه�w�e��z��c���_���kx{���������-�m}�����S~1<R^�=7�����i|~o�w��I��llx���;�>i=��#û�%�c�������S��>�/�?�R~��W�a��W]>�~��o��=7{��f���)��g�_�O�w�!�_S�u���*�W���q)~M~�GZ?�>��y�g�')��[?�ߺxH���ku}��[���i~M맔oW�����_��Ew=���{����n����R���]y��ߴ����=9_O�os�����v�_Ɨ]���f��h���̟�~j���?���t�����M�oR���a�>M������~t��~`ڏK���W^�����oxJ�Y��)?t����,����~�>��o�H��i}k�Ay�zxu}���~cu}N���y���~�O�C����ۿ=��)���b��/��!�ߤ�%�����z�'��i�t�#�L����]�|'���H�n��k�~q��N����Gʗ�ǫ��5�7���G�?�e���ٛ�J�֕�{� �o�������K�W���|��Z��:�/V�����`���X}>�֧]�N���7Z��������K�n=�=o�懴~��o��H�}v��*뷬>���)_����C{p��V�c�Ϟ���������=_�֛i���3�'������긾���O���d��t����?m�9��������������L�i�������_����S��=���Ki��~���OϯV�3�|e���i~4�8���w�/-�/]����n7���ӭϺ�����{�w�y��~I����|��?M������3�?�����i<�'=���oi}`��������0T�W�i���Ǧ�N�߽O����H�ѭ����R{���n?hu�-����I�O���������Ư)�����|���O�~���~��o�����I��ymʧ����׺�E)����q����ic�Ǵ����yO�?�'t��'�mc��?�W��I��n�>�/�OR���0����o��:�>?�x4��}�?��œ�S��L��S�u�3�?�����a�ⱛO�|�֏�'��*����K������W���|a�_�?������W�;?<�<'��Q�n5�ϫ���u���M�t?N���UZ�����H���_����z*�K�����4�w��-^S�M��ݿt�)�w���|�����i*ݯ���n=b���i=��;����-)��c���ևi}��y���ߦ���k�yV䇴�b���c�����.,�����GR��yS���c�|��7��.����?�w�R�,>S>3{�����?�G���Ӿg�����2?��7�b�C�}o�q��)�˰7�6?�7{�s�kc[���=߿��Y�A{�}R�zS�_�-�9���S�S�?��d�a�y���������&/�'6�O�/�S��?�Ο���[����~���k�[~��F|�U[�����.�~,�o��GyR�3�,�-?���4�Um����!�)v�ox5���[Z�Z~I�����C�o�k����1׳���cެ�I����5��T_��T�S������!����x7��_R�5Y}��C�������5���|��'�W�^3{u�����h�t�i�I�Aƿ�����O�#ţ��?�/�|i���/�7����Qu\����_��O)^������"�/�W/f�n�)ݿv��f?�'|��;�˴���J����$���|��o��ś���K���3���-[}���L�����?�߭��kx����R�_R�K��c���t����|,=��֫���y������ö~z���3��iϴ^N�i�w�_���=�=�~q�?�O��̞��i}e�����Q�Wi?���z���)�O����)�?�Sʯ�o�f���ix����O��M��O��Oi<w�c�~y��H����7�Vߙ�������,��?��9�wu����ꝏ��Wڿ������yq�ߵ���4���k����;�M����4_�������?���;|��V������U����c��?c�������ߔ���)=�K�/V���閯R��~���J{��W3|����>b��N��������4�WǛݗ�z6���޷��U����z%=_3�O��i�e���m=�_�g�~��y�H��t�������ԧ����������������t?l��=���*�ov^n�0�K�E�'��4����'��t�/�xNσ�į�k�oL��t��7�z���Rw뻳�[��1v����~,��W�74���z������v�e���o���n?��'�W�~��c�|�޿��t���7��u�������a�@����7�� �����R��o�`���x3>�:�������-��ɗ֣i���oR�����O֯M�A���n���4��x���~���J��+���&o�>��'I�W���~E��M�7��C�/=�0��|5�O��_�ߴ���S�3�O�+̾i�����;���e�7��5~�޷J�OP���M����a�2���2���~YگN��w��V�q�$���|��U��Gʷ�g�'�/����+������n����֧����t}�7��랷u����y�?�z;�c��Jz?���������?�xO��-�R<����Z��ܴ?�����g�^Z�Y� ��b�l���:�����O�i�~��3���A�'���Qf�?�֧��eʟ��}��<�;_�1_��?�y����¾���}E�˴^��g���H�#�i=i��4��R>�:����ԵG�����|����'��yDz^f���/�?)��O�|��4�w�����'=/��w����UY~�xJ�5~����ߥ������m?\��7�K��i<����')�����Oz_'���)��Lߴ?oxN�q)~-?[|������)_��%R�N�ݶ^*o�?H�-=�ZݯH���~Y���n�N������k�Ӵo���n�l����[O����}�����C�����g���b�Ϡ���R~�}8�����������i��7��O�o��˰�k�������ϸ�$����ܑ~&/�����6?���|��pL{�����q*�a��߶>�s�����7�s|��}�-�,^��]������o��Sj�.?r~�?�\��3^)��k��v����Ư���aߓ�S��������kx����m~��&���w�?��L�(�G����c��0�Um���)����]Z��D�϶��#�/�'V��I�=7�ώG~_�Ż�g�H�G���o�w�w)ߛ�����oc��t?i�����i=ۭ�l>�'i=��/-޺������U�������5�5�������g�7���4��]�~��uZ��O��ߺ��g��3�{�q����O��)_�~O]y���.�oY���sʯ�|�龜�/,ߦ��t?j�f�t���7|�|�龜�����ZZ�?������ꟴ�|]~H���yRZ����������������O��n�J��|.�t��e��ô�e��t��z�֏i���#��@�O����+�����֫��~Zz^��Sl=�k��i����4�R{����y��4?�=��f���#i=��w���m�d�1�w�����/��@��yw�~w��Η~߽��=/�פ�U�n�����c�<-��v���,^�5���v�j�������%��W��-�e���+�/���V���)>�z8�o�)_�����"���[9����?����n�#��v�!��Kʯ��^�/O��i�qu�?�G��	)^�_�����4~M��>bZ��������>O�/��Y����,�������ތ��~��?�?v�)_��K담�N�7��)�;=oN뛴����:�W�k��YS��~fz~a��K������W�O����|��'�O����?��-�R~�x��˻�W��?e�q���?�/����'���7���NڟI��i|��+�G������3��l�����o0~7���+�ߤ����|���~t��K��t����|ec��v�3�O/v>�������l��_��k����N���L�����7���n>���J����ߧ�e~���w���^z?�k�g�^zޔ��������K�����o|�����OR��~p�l�exI��4��^V����t��=�����i��ͧ�������t�m��|���?]{�����������~ ׷�0~J�]z��ϫ����w��RZϧ����O�'��7S>��M�g�?�~�?ӏ��m�?�O�|��_������k�OK�Ǥ��k��H�2�O��פ�L����t?m�����4>J�˻�x��I�AZ�����Ϧ�Y�g���<��i��o���I�n?������q�H���&��Z<��=��{L^�/;�����[x>��_������[�\���,�+������j�����	��|�>�����|f��o�U���\����ԏ��}���_�}~�o��䭃��~���s�;�>]�c�O�?ǆ��=i/��C����5���6�>���Ey��7�S�&?�ύ��>�7yS|R^�+�������yՖ���7�S�&_���,�S��Z�K���}ʿ���{�3�-�ml�j��Y�fO����{�/���/�'�>�|�1�a���h���~)X<���e|i�Q�߆�oƗ)�t���G�R�������x4�������x2�����S{������)�=�����i���i�g�3�g�o�O�Qi}��EZOZ>����g�o��,�p~~��m��V_�����;����g���t?��k�'柴e��t�d��z/��X?��w�'Z���������o�A���_g�2�4������������ݝ��צ����jx�<�'�Ϥ���g���%㷴���w��o����W��5�����U����ѭ����ɟ�o���勔o���� ݿ��U��w��Qڿ0|_�>�/�;H��)�-������Iϯ-^������S�Y??��m��-����t?������t����z��'�_Ƈ����}���~��Iʷ�?O���߳~��W��M����3�_���i/�?����X�o2���~*�������`Z����,~�|�����'��}��U�3����_Z�H���~��C��Ç՗�����֟N�oZ�����O�hύ_���7�>����͟)�������d�4�ϥ��X/v��h�n}��g�����I��i�$��a�k���f��<��3���֋�O�������e���*�wV�����?L���w:�'oZ�^��4��0ۿ��#=���HZ_���{�0��٭?���S>��W�{�t�;Z�����c��΃�~Cz��;폦�����K*��#=�L���-����xL�g���u�ä�]�R���B�W����^N��t?��GM�ǥ���j�L��i>I�%i~O�c�]>I���yG��V�u��Sz>`��t����M�Ə�/1�������N��s���]z~���R�Y?��qZ���Q6?��E��������?��t�����f�t���K��jz�D>�xL��i<Z?$���������W����翩���Mi�����~@���������/�����/g<��=��;=��Y|w�;��ho�Ϧ����_U[�Z>I�t���i=L{��״2{_�}ϴ~M�s�_�_�z*��ؽ�g��z-�'���l���;��`�ף��_I�~����{�S��~���gu�w��ez�&͏Vo3~�E����C��~���V�>��M���l�?4{�|Ʒ�~���������=�i��o�z�?׷�zʿ�/��e�}�#�_��K��M��7+λ^�����O�o�oG����v�����5�o����k����#y�/����I����Ǿ����s��s}Ë�Gy�}������Ɵ�����9�Ń�gxH�O�ͱ����|nx���d�g��������6�o�X�0��z/Ծ>J�œ��3<rL�M�?���{���[<Z|��%͟�߆��f?�����M��#�i�h�H�f�Ə��)�r=�#�wZ��|`��w����~�䡿�|g���7��ċ�o�^R�X������m�}Z/���n�N�����K�2�L�h��4���e{�j�_H��/i=��o�}�?4{[���g�t�e�������i~���~���1X�1���_Y�����&��C�_�\=N��S��t?��Si5�/ڋ�~M��޲��{���[R>c��|��&/�U������S����c�'i�c�O^�i���O�o��������4�/��i=���ɴ>6}��b꟔���C÷���#֟'���>=���+�o��~���i�4ߧ���4>6>L�+�<=��,���~-=�����'U���n�'�G��,���ӧ{��Ώ�����Nϻ_Ə��}o�랷����7��?�}���/���׭��4~K�_?���ݧ���8����8�/����g��L�?���=_������c�5����?l?n�K�?��)i�3=o�:���z��`x��?���'�^�}��'�'���'�����m�[}^hx��v���Ou����S�~3�O�y�~!�'��m�Oz���|�}��}�C;�ꞟt�S����ۭ��|M{�X}����L�7���4�t������o�~�{�h�g���w�I���GV��g������=?�z.��[�4=?J�#������iZ�Z�I�U����?t�Y|w���Hy�����UY|�����?����������'L￥�gÛ���U�Gz�"=H��{?+���/���|�֣���}��5y�t|V���v���o��==����N�)�Ǵ^7�,?��'���|��K��)�Z>O�w��Ezޔ����+������c�K��Vo�|���Vϥ����"�_z���������|���k��gf/���?����}��}�4_u�����>��;���k�Z2�g�?3���E-_�~��Iz�b�W�ݯ��6�7���nz�G<�yAz߲���GY|��)��iߴ�J��?���~��������||n�~�׫����:���ߨ}����B�����~���>`�%_ѿ�3��Ń�۵�7�5{�||N{��l>~o���9?����������^|��Q����1�y���=A���^�Ԟ_�G�P���wϞվ�o�g��������|��=7{�������e������)��\�����������c���-p>��-_�}��-ލ��9�3p}�#��1�3>��1�J�1�k�����3�����1<Y�`� �����ƛ���������v�<)��}�y��������3�/V���BW^�ߔ����}߭R~����;�/��7����O��ݻ�ɛ�'�����������������W?ۯ���4�}��-�>ǆg�͞6��c�0<X�g|j�|�Ƕ���b|A~�s��4_��w�����~�L����t���h���i�5�o����c��?J�7������ކ�4>�/M���o[����m�1~2Y�ӟė�?�o�#���O���Oϣ,?0�sL����g��Nj�W�c�;�7|X�j���<�����i?�ۯ�?����������3���Q�4�X|�>�~Ϟ�����Ԟi����/�}�����Z���q����������L�g�E��J��fï��m?`��/�}l�����'[=k��Կ��wz��{�����֯J�A��~��w��f����D\��C��V�Z?����d�Mϓ�d}V{��o��n�H﫥�~����޷~��c�3�����3��V�[����y"���������_�7��������S��_l��������o�����7��gR�����<!��)���z���V������Z��ξ�������6��S{��������������~V���)?��'�������'�߳�=���]���N�I��i=`����|���z*=OI�t�{-_��)���c���w�m��򟝟X<�-�������ɓ��;������~�͟��ߓ���_ꛞg��?��Z��~)�����?���Y�]�_��V��)�}z�g�����>����S��5�����߬���^��2{�����;,>���4X���&��b|n���쾕�g�`��������i�f�1����2{Y<X�N�#�ߧ�~ʗ�}����Wv����h��6>M�Y>��T���>�������z���������>����[�b�Z���O�o���n���U�?��O��J�O��wV�y7�t�o����N�g�/��d���Vߤ��]����i}��~&�����W���Ez'ů�Xo������f��x��2��O����i$=oN���^��2y�_h���޿�����go֞ψO��Ń�9~�\��~�>�=^ٟ���P~�o�߽s���~*���������z���%�X?0���M^����>���>7�p=���;������A�Ϳ������k�ml�7�������o��i�"��>�7},l>>�=���������'����ߌ��|~'�}�����8?��\���|o���o�j��������},�_Y�`�����W�/�o�4>��i|l�0>��i�u���'{n��z���=(����N�g���������%śŇ�i��Vo�|�������c��Cf�O���o��Z}��{�n<������e��/���Y��|g�	�G��-~�����>�/��z��!����|��+l�a�Bն?űً�M�a�[<[|sL�Y}n�J���=)�̞&��ZoX<S~�o�-œ��z��e�1<������;����K�g�7�����+V?��yZ/u�/V�v��i��j��_��-����|�o�x1|Y|��)^�����ջ����1��lr���R{n�S�'�b|b�Ѵ_e����̞)_ߧ�n�H����-��7[/�WV�Z|Vm�����y����t�"_�~&�o�������P�G���k�Cz���m�1y-��y��#�Ay������~�=7�K�)�7{�?��g�-����R>���B��L��&_����s�Ǵ������ꯪ-~v>G�8���>i���{���I�y�����Ɵ���#��L��V����~�ٛ��~��a�e)���5����;o���7���~����Wʧ)�?w�۳�?��7��O�\?���������_����U�7�o&o�>|�/L�z>�v��{��_?�}�����R����o�gʗ�Η�/I����~��n?3=�$���W��v�n��{ó�գVO��{(��t��=��:>�z���������8�������+����Xz���g�[<���~��;=�J�;�~�oH�˚>/U���O������w�~$ݟu���������<��ў_��Z�G���ޏ�����������H�����M������vg���#�_����+�7��j�g�f���ǚ}������4���װx�:槴�d������϶�1y�>Pz���~�Y��O��~"?s�L��>���z����߯��ߟ9��������'�����?�/�ק������\�����rL}�=�S~��������rLP�����?|��8��O�������χG���f?�o���3�z�����3���3��o�Ӈ��s�o�OÛ����뉌��˿�=��?�K�k�l�������.�+�&^��ٗ��>�k�c�6~6��}-�Y>N�]��V��?8_�6��~VY�m�-�?f/����J��{��������?�?�'�����j�8���M>�֋��g�ex����OV��P~���_,�-��/�����wϞU�j�o�z5�wģ���7�_���1?��|N���_�_����l��������8���_~o�������K󟍍/�/������?f�F�5��m�o�[[��_i�0<_[��>�7��)�?�/(�����o���3Vߘ=�~N�#�|i�e���i� �W�z?��~i�����i���M�4�X�!�u�;Mߴ���m��������,?�������k|gx���>~�����ﹾ��[>K�����w��n=k�
ӏ��>��O����&�ŗ��\����+�?�O�?,,�����w��i������Ϳ�����1�3���$�ô�ʿ�~zz~lx����w1��ߍ������&��+�7������^�������Z����J��i=a�i|yg�g�/�5<��`�7|Tm�������v^�����Y�/Y~���f=e��������?�?���;/���x�|���V��8���y�Ň�Ӷ�3�t�����mb�9;�5~3>0~��D���������]��o�-켁�s�w�߬�`��忴��g����w������������0������+�����>��Cz�����$V��o,����4������,��;϶���v7����6��g�6��b�����9���6�=��������m>��n���d���O�'�����OZߦ�����Q��������H�W?��%��p&z����o�״���ƻ��^��|������Vvޖ��~S�O����VX������a?0=�2�w���a����6�=~�_�z����-�o�b����|����|���M�ש<�_���o�G�o���O�?׳�4>�=�f�����Ǵ�9V=��\�}n�b���߂<w�����0߳�b>!?����������������Z��!����|�������g��7���������h=���i�s��'kާ�y�����{�������A�s=��1^�������<\��c���\��Q^���e����^ԏ������k|b���Ϝ?�k�O<�|o|L���1}���ɛƧ������9��c��s���f|Ay,�?�<&���VX��|Ƨ�O�9�a�����#Ǵ�c�G}^�����n��?�ʏ������s�O�q=�7���ɗ�MZ�|&��tc�d��|�1����������[��Z��86~�xM�3��K�g���)R�t?l|��f�����{���^1��|��f/��x�zؾ�|��N��|����s�_Z?����}���I�_���ύ�|O�[��}Ο�?�����?�������7>���KU���ϱՃ����`���^"��	�7�?�Z�J�R�'�=m}��������|����C�o�m���V_���O�>��s�_�|����|N�����j|L���>뿤��ql|��猏�<��2<_?q>�o��8?�O�i�+�˿fo�k�Ӿ���7�S��&�������ה���7|s}���Oyȟ)Y������H�Uֿ1��ߍ�L_����nz�����~�ū��쓞�v�5�Z�l���ǌ7�s=Η�J��i�����_���~DՖ�S�q}�ϔ�����Oy�|�{�h����N�g�3��S���g�2���Vo���'����I����֯5�t�;,>���`��|�}/�4���4~��Ç}߽�d���m���/M�_s�4s>;K�-&_z��ާ��7N�u�Y�o��|��EÏ�3;O�z�_z�<��k�G�N���zvݵ��O},�����_V?�?�?i���r>����ָo=�m\u\�����+�oX�`�<��X�.��g������y"�m�Y�'���U��k��{�����gύ�<!�����~�K���}�OZ/v�c��su���2����l��<$�/Y�m�����F{Y��%VϘ�i}��������o�����"�_d����>�󧝷��k����Sz���+��{�����?�~VO�y2���v_��Wն�2y�^O��8����o�)����|@����!~^<�����W�ϛ������߂=�����O~�塼ԇ�S{��~�H�O{����Q��~|���>�������y�����q~����/�`�����c[�������}����|��f���8&���������||�����O�����#��e|��o��zm�����������������|j�����1��3������[��'�/�'�g��O��M��ø�`��Gԏ�4��_�o~����[~1����>�����?��p����x�x��Ư���i�n���0�?��q|Q_���=�o�菴>4�������l����/~��M_������c|e|d��M���V/�����#>���G�Su��~����V_��\�η����������k�_4~�x�|a�`|`�d��9�K�I���o�?M���>�s�7�G1>������J�3�o���6���}���`��:ޟY<�}RR�_-��GV����O�&���,��<�����������=���cxO�ħ��;O��-����_���|��[�sl�b�5�?i?��X�J�����~����m�b������a���_�߆�?��^�_-��H;�����ϩ�.=�|_䫪m�e�<�����?�?�x�z���姴�o�f_�Y<[���ޭ�H�K���3,�����O�Gp>���2>�f�����c���w���1�/��2\��{���O4{����o��?G��y`�_L�o��Ξ���Ń���ޏ������|���OzQu�?2��~��o�7����\/�������S^�����#����_*����_V_Z�!���~���5�פ����ްz��A[�o�ߔ��Y=g�����=�~��׭��|`� �O� �����8�����V������b�?�����-�Y<�}|ç�Ky����v? �O����˟�O(������j���i>���~����>@�4��������~����S�[>�x��j�߷���c�Q>�'����?^�ǖ�l=�-�޺���Cz�g�������c�?������?�������~��[�����[���o��z����}T������}˧�_��H6����~�Ջv>�z��L{ql�oi=K���3��Ʒ��'�O���=E��[������@~>�x��xc=@{����=�=���7�&_p?���c�gߛ��������_���]����?8?�g�P�C�8?�'k<+(ǜ�c�˱����&?ǯ�~�� �-��G�������\�f��Y�������?��c~o���)ǌ?�������[<s}���i���6{X|�{���g�s=ç�9�},r>����x3}���OV������|b�0�#�9������i����a������R����g�ǌ��>��K�	�3>�z������I��<�G�W�|��g�����ك�������3�_��<V/��4�^�m�����/���ԗ�R?�9�~��o��Շf�??[}����S�W�\��u�c�[�nc˿V�Z~�z;����>���!������Ϫm=��ϖ_�z������/�~�߲�9?�A��|l��埴^b~���7����o\��O���}�ճ���>�x��i��V/Y>���+��pl�5幓�Y���,�p}�������׷�f�a��Ə�W�����g�����|��v>d���o���\��m���/�o-�r=������~�_I�g������<����M�����vf�[�F�86�����s;����O�����|V��R�����1߯��>�������J�-����&��yw>���F��=���������o�O����S~;_�xI�7��?]{Y�Z?(ͷ��V�3�h������[�H�ˬ_���Q����wi>g=��w�<i?5���ݝ�R{����ű���i����������K��Ɵi|ql��՜���Ư��N����l�����^�y壽͞V�Q�O��n��{_����o��8=���\��:���|�x�~��4�Y~�>i=f��cZ?��{�ǝ�Gz���W��@��S��>����oV�Y=��������o|`���S��sL���m|g�5������l�c�g��C��-��Y���#�>֬���W�ȟ��y|g���?�}}�z����t�����j�?��=�Ӽ>�����ֿ��C����r��?������=壿�=塽8����l|���G����~�hO�K�9?��Jm㿞����7|p}ڟ뙽���뛽�>xN{�f���s}�O}������i����w�ó�KY~z���~�u�X��v�O���1��|�?���-���L~[��[<Y�q>��#��}�GS?�-�q=�����^&�~�W���/���8?�s>�����ҾU��E�s~�g��o|@�-??������������a|��-��=�i|g�I��~����[�t��M�w�69?����6|�<6�E{P{N��x7~���>�X�o�M����z����Y�l����c˧�'����g-�����c�'�m� ����o����磿���{�O��K�)��/�����������C|r~�_�^�6V���޳~�Ư�����ؾO�qS��s[���|�G��s��2�,>8�~���1{���������������fO~���3����G�c�o���3��1���)[~�?�Y�W���d���G�'��}��ix�:��|n�?���K{����7�����k􇝧�������Oy�7�H�7|����4Z}M{Z�[��<������}h;�H�3�>��+=�~��M�������>����c���pL���y�������V�Z�6����Ijo�����Ǎ?S�Y=n��T~�3=/K߷z��������\�·���N���!�~�~�ً��}��?������g�O�V��ؘ�u�9�����%���߸�����{�#=O`���i�m�֟�z��3����Gz?����M?�����2ۯ[}�1�c��ƣ��i����K�K���N�Q���Vj/��/�������J�C���<���~Gz�,����v����~��_�o�����?O���ϖϸ�?V�����>���>|N>0i}���>�C}�<���c�Ծ>��{�}�ߠ��W�Y��b��w�p�s��������_?8�����W���z���#�����~o��Y���)/����=�������'��<|ncڃ�>�����R�Z<Tm������O�(��g�3����۞sL��?���_�}�}��5�q|�����z�?�|���g���ă��1y/�ǜ��5�q}����>���(��k�I�a���5Q�g�G��-?2�9������Ɵ��^����_X>���Ծ�w�'��q�'\��j����=��">R~0��>�����f������oϊg�?�n�_��ٓ�[~b|��>�g��B��ǎ�C~��V��~����A����\�����g����c�k������W�φϛ:�����O����wڟ듏�hO�_��s���|N�Y|Z<���)_/VoX���B����/ڛ�?,_�?���'���9��x#��f�7ˇ/�����_e��tc�3��:�o�O�����|e�A��_f�m���L>�;������q?e|o�?���/��O�Y�Oӏ��|`�a�O��������կfO~o�e��s��/�C�_������?\/=�1<X=��k���7ϊ���������'�'�>�%�h��k��y��/��t?�=�0>���y�O���k�N�)i������z�����Vߤ�C{Y$ݿi=���/�� {N}�^Z_�s=�'��i?�����}z� ������x���_����V?�y��'�~�z)���{��7y,�1�}��m���m�g������ݗ���Ova�c��z����f�;�Oԏ�����=�|��X������)��ω/��_���O�76���|�c������O����c�3�K�o1��~��;׷�|��Y?���3��}I;�5|��8�a����f�?��H|X}a�'��1���8���[�rl�?;��3�/�_�x��[{>����<~�����s?M�1�o����ȧ�G�����F��=�y>ڋ��s��甏�ў�ֶF��{��Zm�������7ǜ��p~����/��f��=���sL�qL���|��ڟG�x�=9�a������%��[���z�������}��J{�{���s�Oyh�O��_?��,>(�˵��w~�甇��_���d�����k�I�>ԟ��|�'�כ�ׇG���s>���q'�ƃ����O�1��=(�����|m�����7��W��oÛ����^�|�6�}�x�x�z|n���a�'�}��(�ՋO�>�[���R۟��k�!���[��~����į��������9��C6���߶����o�����i���w�-��	�׶?�}��0��z�?�K��^6���/�1}������7쟘}�����D{P~Ã��_`�h��Jmϗ�ll�m�g/|N�������b�D|S~�G�O�~����<�5�[���M>���������|��R~��o�����z��}�m?g�Q>Ƈ�si��|��?,>�����ٗ�|l��~i~���'~�ʓƏ�w��)�S���Ã�8?�z����Y���������[~oc��YO__���M������������+׳~����wگ6��?Y}�������{U[�I���az���(�I���n�?��J����s���N�g�'V�[��������x�~���h/�o�����|o�r~���7���/�?Vǻ�[?������;��a��������3ԟ���9�z��?�ϱ�9���^���y��;߷|a|����}Z�p=���/i�j�]z�.�g����Y��c��,�_�U���'����x�},�Z?������X/Y�F�Y������{֯���+=�z|��O��A����g�?b�������S����_v���|d�3������V����������4��N�Y~ڋ�A�#x��Ń�����z����W{~!�g>��)������J{�6���ԗ�����?�=�'2�g?ڗ�����F<1?��c����l���П�>\���_�|���o��������|���~�߾�z���F�x���o��ƿ�W�/�k�`��zď�o�'��~ox��f�9�ٗ�������?�W����o�HZ�?Y��s���3{��-�9�����Ɵ��i�r}��h_�cx�s����4ޭ^1<q~���+����׷z���?ă=7<�~�,�m�z���������8?���%�_�gx����;����>�_q�te��|��-_П���3��߰�����s�����q�W����O|n��P���Q��c��a<?�{ƫ�'��|�և�/�~���_����j��'���0���5���/�w�2Z=��!���7u�w���d�7����`c��X�f�j�4|����ԏ�о\��ڟ��%�|��g���4�{ڃ�3�����o������<����|c�e��[�Y���O�/������#���k|G�Y?��Mz����|�ϱx4|[?����{��=�GVp}�O̟���O{>���z��퇬�a��4_�~��@{�i�j���h֗�{7���(��_��������`<���,ߐ/h��:�������ħ����<�g�f���'��g�o�t;_0�Q�������OƧ���[���C��<��o[=h����oz���?�'�_�}�o�T�/��l����7��>�|���k�ߝ��������#��z���7�������	쿱��9���3��7��G��=�w���^"�����ɗj���������O�c���9�G{R~�Gyio�k��<�'�o����>�|��Qڋ�&?�_�ֶ����?R�������Oyw��S�Ǧ�{��������'��?L~�7����������>f�o|d�S~�K�P?���?ī�����Sڏc���(��q~ڟ�1�-����ql�k�p��;����j[1�S���f�g�����9�I����+����[�����/�1Ӿ\�x������n������oL��c��o�=�b�����3�c�9ף��?�o��;�����Wu����?����3~�oh/~o�h���̯���Y��x�x���>�1�7~3��O�9ף}m=�3֯���ŋ�iO���[���i/��G�=���������)��o֟#��9��ǖ�i?����O���������X=���t�`���1{P�����K�������o�?Ɵ��|ԟ������;Vrl�-���G�S���Q�w>��|���)/��x�|���}�/~o�����_�����O�3~O��}���������Sӗ�a�����?V��};�����ً�X?���tb���K���O�G�r}���:ŏ}o�����1����������6�~�Ϡ���K�!�c�0�>���oY��z�����~[z�o����G<��c���~��)Ɨ��%����9��k�=��0>�o���|�/�w�'=O�l���o�CV_[�S���Q���ǖ/��+�?J�{�������U�������v>c����Gz�z��A����~�����ԗ�f�^ma�y֟�z�s����h�������w|N�z�����B�`�e��v4�GЗ�q�a���������"~�����}��+�?od����{[������9����=��f��:�۷�����G���������'ק����R��>������ڞ�Tm���9?��?����B��{��>d���9�?|?�+�����?��O���}~8���R�_wĿ��O��=�a����e�c����zo�~�}�������>�Ay�G˿�ק~����hO�/�1�����;���_����?,�����->���7�a����o���;������s}�|`�g�R�o�o���|���z���{������m�}S����/L>��|B�_���7��cï�ϩ�����z�Ozdoÿ�C��޲|tS��)G�߷����|��c���?�����߶���ĳ�ۖ����7L^�����h�0�Ҟ�~�����ŷ�'m�g����~���[�?�o���S�G�?�/����c�w��>�x����Ϭ?g����J�M��V�Z�M�����<�w��Mm�L�H�1�w��_�׳z���=Ƕ��|�g�=�<����ӟx�z��w�/���m���ԏ�����C��96�X?��#\�������M���:�>��������i�����/��)�7{X�����q�}S���y}�g-^Ɵo�o��3>���}���~����o|�����t�d�I�{��[|�Z}M|X?��b�P�?���I[/�'����O�ߖ���c~JϏmj�$[����K�o���-�����ߧ�ƿ��m���3�i����]ß����g�wf?���K)_��@z�g�M�w>��a��`ϛ���s3_]f�}�?�}����|A�|�`���%���9����}ڏ�i�?��z���K���8��÷���B~���|��������j�{���H}�����z���sL��Y��(<a=����ě���}��M�K{R�����߸���x"����/���-���c�c�k��jm�_�S~�}(/��)�#�=����hO���?h��;�x�|�x��I<��>�_�7��P�~���g����'^�o�S���+�ݏ�ԯ��}o���`<Z��F�������<����g�c��s�C���(�M���/)������-?r������M��{T�����G��ާ~������ڃ��>�����|�O�>g<�����x����o�������V�����|��K�C�~�^7u���s���_������瓃�|n���?�A�����a��{�Wi��c��_���='�l�m��K��}�+�����9��o긟��Ɵ��j۟�~���;��0�5>%~���,�����6~�����}�o�׍����z���ɿ�'�����~2�o�3���s>��Z�����nxL���a�XûՇ�/�3ף>V��l?b�}����-����Ǵ�f���	�?�����������_7��>|N����i_��4�m�6����ws��������T������e�?���P�����Qi�����>����~��cۿX��|l������~������V/R_�GV���<��k���C�'�o��M���,~mL��=�?�M^�_�Gv^��g��2<Z���3^i�g������b��'��l?b|���9��f�g�/�c������ۏ��f������v��͏�_����\�?v���e���[=c�}���c���c��b�R���i��h����;�z����߃=����?x�?��x�q��'���y~���S����f��9<�g>��6�����Q{<�������sڇ��z�>�C}8�|\��|�'�i�/�b���Wk��%�@<^S�sL{�|��?������~�/ڏc�Oy�|�������/��1�k|ʱ����g�{�|B{��>�/�a�>��\��Hym=�O}(��;�������I}h�������}���#~5>���Զ�`���o���->-��>�姿(�)����x������-�2~)�7<1����<�g��7磽�V�x6���,��?����k���/���'^h�k��<���?�WZ��~V_����[���|��6y��,����O,��?�'8?�E��_V���V/R>�	�����mF�io�_��7~o�����?�G����������}�o����%����z������,��^H���/���c���|e�Um�-�g�CZߘ�������s�����>�_�=���~��k�w��e���j�G�W���!�O���ڞQ��-���������q�_3�1>�~:�m���whO�S�W�'=H�i���h;����/��׍_(��o��w���[=e��t?f���G��^\��o|i�L߿��>�_�7�uS��v~?����b�2[=E{s=����\��m�/��ho���9�����'������d��O�_��R_�6?���|��𕞗�~�ϭ��v��q�G~L�#9��U�z��I�����3���Y=f�i����_o�Ư����$��X=@��~������v�����oa��<j���e����w��߫}�&�s�K��������������;s|�<����Y�O��O`<���a��c������8�+���a����>o�����)Y�?����K7�������7�r>ڏ������������u���>o��|�Ń�i/�O�R>����=(?�d�S^ӗ�ioӟ�hSӏ��}h_��=��4{����ߟ�|F����f�C{2��/����K|��-���m��1����ԟ�����m���XOߛ������V�q}����|o�Z~��-�������Gړ�6>2��?�?�M���>K�����5{2�G��/��'^��ԇ��|h�&��z������A�����#3�R�o���S�����L��pLy�>�|b|b����VOX<���c��k|���>������8�A|�{���:�О�֯�}̿\��f��|h�6<X=a�h=�ٳ�)ǖ������������J���7ߧ?,��-?��I�G>�|������ڏ|�����3|?�~�ڞG��O�?�z��-׷x'ߧ�>�|�Ǵ������A������S,�������ǌ��-߳?M���ճ֏��L����M{X�d��~��;�K�{�/���9�a���Y=m|xS��Z~O{�ԏ�Q�S��[=m�����=���7~$����������o���uz�h�e�w8�է�o�_�S>�ǟ9�hO���������E~����g��k�S�;���_���	�߱~Ez>n�n�-�o�~��_�/�o[}a�6|?R?>���w�����>E�Y�o�>3���3�߯}}�z�������߬O?8�/]�����f{�T�x�n������?�g���3�|:����_ڃ��9��񛵯�_�'���r��<i�p}����K����{��x����cڇ��|�3ǔ���}���G������|L�����|n���o|N{r��oj_o3�|O<s��h?���O������7�Q>�'Ɠ�?�c����c����>�}hڛ���fo�cx�����4������Ϝ��Q~�g���V�ѾoԶ�g|F�����iO>�~\/�;�G������|6?�>���|i�����"����}���,_����-�8N�iʗ�#�m���V/����z|��Q���}���_��VS_ڳj�����Ǿ�=����ԏ��|g�f�iʗ�_�Cڇ���,��������k|G��R�'m�t�L�,�?����g��x������0>��7�3��P�����r��9���3|X��~��|f��O�~����/�o�g�������/���|��uӏ�i?ۿp=ۏ��ߵz��R�ߋ�o�������|�?��v�@���^V/Y����o�`|e��ŏ��c�q�'�{�o��������������	�3�3^����֏��#�3���������g���	��?�w;�H�'��/l�����O�g֓��sA<X<?�yz~`��˱�o�hZO�y������>��=�'�CyiO�G��<U������+��`�/�'�f��?�s���xg~����k���c�I��}Z�a}�x#�S�+��y��z��j�d�C�1>��G�s��?�П7�x`��F<�����>})�����3��3�|��G�8���s�?�����٘�����<�{��}cڗ��}��1��=�}�����L^��Bm��x����|������=��7ף>�������+���9�J�h/�?��������S>~o|c���P^�;�7�2���_��~��S�7k[oƏ�'�K��Z�������y����G�d��c�o���������':��>�O�^��˵?:��8?��<�;���l~����zV�ў���|�O�/,2���'_���^��m�Y�G{�����b���1�3>y�������ﴏ��������z���|C��1�[������Ə3~\�����7ۯp=��'���~���VO����;��z������ڞ�S_���a|i�C�������m�t?g�e��k�0>���7�7��5>b�0��|d|j�1}�o�oj��������G��ճ��|K�s�Gy�z��������6_����fo�'�'�m�鴟C�l>�g���_�όW�G����Y���K|R��>�z��A��޲���O��������i}���C֟'Z��/-������	Η�1Ƕ_5�I�W�_�z�ϭ?a�ei?��xS�x��)~��]�Ƕ"�϶~�?���g}��ˌ���{���ͭ^�z���������io;O"?/ԏ��qw�4�|v��7`�o�~=��{O��'>�߷�9�����ӣ��m��k�������s���Kf����<Od�G�l�?8�_�m|ў|�����oӇ�3�F������ɚ����9?��������|nc�o�3����ԏ�j�O6���g��3�c���io�����oj����?��������a�r��j���/�K�(/�S~�����ofo����S�-�A��}�;��/�g���(���S?>7����/��x�9��ϱ�������h�'����������g���x"?������7Ǧ/���3^9����o����|ďՓ�>���������]��n���By�?�\��%�r�b�;�ӿ��E����o�w�_�k���壾7���I�W���O�*����?������������3>7<���ߧ|�o���g��R�����'�mB������c���G~��Ƨ�������1�m��[|[�G}��3}�����E����������V?X�K�X�`��s�o���ߛ:�'������k{?�����~��5�H�a>�<w��{�7���O��j����͞�'V?Q_�Ϭ�d��������� ^�����c�������q>��p�O&��7~�����x��V��sƯ�o����߶�6/֟�z�x0��>�?������h�Sʟ�W����{������K����o��t��M���S��>��t�g����7�?����ğ�W���?�/�a�e���n�շj�"��o�g�ǙOy���5��3>��~a�����߬m��q=��R��}�#{��~R�~ �#���ά��+�9�}�g���"�o��k��+����זo�__���{�K{�^�_~��9߫���C�9��ڛ�9�����^<��cڗ��|�{ڋ����CyƟ�Oふ9?�O�>��>�+�#�i_�'���sڛ�3�ߩ�����9�#>�>���pl�{����w�����K}���/ڃ�0>��\����D��/����Ļ�/�s>�����9�My�'���9�7�ҟ���x������\��4>��/׶>����>�������7�'�>�V�P~��c������GƇ��C}���U�7V>L?�Gy��O�[=��ė�hO~�x���'��|�'�9����ԏ�@yi�G���-�}ڛ��~���c�iO���}�g���_�o-���������s���>�e�`�#�����iO�?,�?��x����i���c�d|�q=ڋ|����ϱ���+�C�)?���i��/�����?��Ʒ�_�/0��^��������������7f_��������M�{ƇՓ�0����|VoX�����8�����cx��6�c�K�����V��>)�9?�k����1�����Q������:�G���K��~��d��x�?��;_����M<?��������g�������7�?�{���^���w�����_�}�K���o��{�� ��_�7�c��������7�����������y���Gb���G<���{��7��x���S8�C��>���z���D{���6s�G�?�a�?�K�i�K{>��m}��>}�������G�L��s����1��=�_�K���Oy�>��s�������D|�>�o���������|n��V���G��1�=)��?�;ʟ�﫵�_8?������=,�Ѿ���z����o����|�'������������{�G�������Ɵ�q=ڗ��|��~?vT�r=��?�ñ�O�_�Ot�oL���8?��x�����}Ƌً�m}�c�Oy�G�w�?��_���5�E{�9�o�������|��ԟ�ҾVo�����~��C����C�6���M���?��i=I��o�ڋ������������W|������s��|�1磿i��(?���%�G�����|�������������z��g�'���O��z������e���Q�7Z�n�G~�}��}�1?Ѿ���$>�a�'~_�����W��-������������=��9?�����?�������3>��X��y�ϧ��ڏ�A|Ҟ��_�×�G}R>������֯��������%�O�ho۟Y?���_�Oa�c�(>7|���?���k�,۟p}��j�����_l���a�v�g�S�h/���#�K��3�ڇ���o����j����e��۵��
��쯲����K�}\����3^�m}�~��g����?���Zm�������_����Q>�OyM~ڋ�Q����|\����ѿ��7��9�=�������7k�u��Jy̿������L_��I��}�O����_����?Q��k��3�����|����ԇ�S?�3�����_�G��>�D�nk������d=:�K�/�j[�Q~��Fm�W�G��Bm�%�#�%ǆ���w��������`>���!�3�h��甏�i?�?b����hO�/�c<p~�Η�����ު�y��;/�����@��ޣ<�W���b����?���1�g~3����~�������=g����Oi�����~��-^)?ߧ>�g|��	�����^��ԇ|��>7����[�Cy�=�����������:�wS_�G���4��{�O��?ɷ�g��������`�������0�%���vi�%�����=�G�O�_1Z?��Y�G��}ڋx�z�����3�I��=�?�o�?���8&��������_c�����)?���i�������W����fO���Q?���?@y�����W�o��ַ���l���2|R^�c���}�~�j�O��������-��}�7�c� ��M_���GV����?�/�v�C������Oj��y5��z������nj��߃8�wk��c�������n'�>M߻Z����g��/����wj_o�~���ב���?����?�����:�C<�m����oڋ�~(ߧ�������/��\�~&����k��C<ӟ�OY�_��?����g��x|�����3�����年�d�b����~?��y}��zm��G���6�h�OQ~�O������7���͞ԏ�ލFl��;��x��ުm�M�mL��>����4�_G�S�����?��o���~O���7��z��+�S?�g���kī��a���G{��ǌ�C{Q?ï�)���c�'�7��h/{Ny��G�q>>���O�3ڗ�n��z�_ڟ��������1�D|�Ƈ��͟V���>|Ҿ���M��� ���ԗ��}���c����O���>�O���_8N��������~����� Q?ۏZ���C��>��ŋ�G���A}����J}�ě�S���+��?>�w�=����/��9��G}����֯�z��E��Nv|���z��-��[���z����M�﬿E��>3>�����x���=߷���Y�o���=����VOZ}b�@y��Ly�O�?���w1u7f��`>��/o'=��/l�E{Z����Q?j���4�����z���>��,��뼯���7�|\��^�����wa�a;�^���y=�C���Y����zh�����އ�<���][|��d=���������}|��s����zT[~x��秔���޴���ȷG��sӗ�E��{������|t0?��<o���W&���;�������rm�_Ӟ��O�P_�'�e��~���P_��1���y��ߞ����s�����<������)�嗑��`=�g��|&/�L�2~���^�Oڃ��|��m>����}������zm�?��%��?��9f��1�3�"~�/�'ho�?���`>Ï��������|~[[�X���{��ߓ�_�/ƧV�S?�m=e�5��W�'��>����?�7�Wڋ���ԏ�n���nk��o���x3��<VoP>�o�����K����ϩ�y���;��nj[O�X�����X}H|p~���s�C{�>�/��zԟ�'��ߓ�h�G������?��o�L��~2|R~�g�:ǖ�������,�����-�h�O���'�9f=f�L�O2>�s�/������37���:����-?Y|����0���о7_����I�o��9����^�_,~9f�q>�_���֯4{q=�q�����j�n��M�s�m�������|߯=~��ǟM�j��!���ş՞�y�|��&��$�kx?�Ń�~��{���7�O��>ߑ}���}�~<���I�)������1��r<7{P�������G�����U�;�����io�Gy�ϻ�����C�<'~hڇ��������兩a�>�_�9�e�iO�)�I�{������oj�Wڟ��_/��~��z���ߚ��+��x0�6���7�3��Vm�a�+Ɠ�����/(�g���?/���Ԝ����_����|�M<P>����O���ڟ���q|r~��T~������O�O���o�sL<p~���1�����䥿�w�G��̟�w�����0{s}�����\�c�o���8��#������������e�y���O������9�E�P^�'��E�/fo�o��c�s>�?�������Wj{��������C�o<����W���X/Y�o��xc���i����=96|X�4ym=�?�n�����ɏ��?M�o�'Qƫ�������me��O}���������K~���G�Tm���Ϗ��j��b=��#�E~��⣃�߭}�J~���nm��<��῏G���X��	���!�-��|��~����am�5bs�k�k��?�W�x�塿��K���+�O���o���g��Z����~�����S_��������)/���{�����\����́_���F����&^���e�����+���5��^������^���$��G��������fO���OtzV�̟���z���9�7��Jm��������|���x�<�����Y|2�����@}���w�G����A��o����=���o�#����_ǟ�O��W(?��p>>����c�3_q>Ə���h�o���z��sL>c<��ԗ�ӟ���ڟ'��S?�c��g��z���?�3~�})?�%~�����s���`�d�$>�?��}���1{o������g�/�'�>����3>��V_�}���ۜ��W�k���C�о|Ny(��'l�k|���������'~�>f�J������=/�~�����eԇ���'�%�O�o�g�������l��� �����K1�(/�'ߥ�Y�_���[��Qm�C��'�e�)��3�Vr=��h�K{Y?��[�H�������͞�8�������#��y�|�|2��)�����~���o��"�r4?�������1�;�~����|�o��;��O�_ڟ�Q�j�߷`~����i�/��x���������zc�/�G�,|~ ?��<ē�c�����>�c�'^�?�����g�g��_#����#vf~�io��������{S��"�#�/��nm�i�/��|�?S?��1�ߏ���hx�}(���o��#�P����>���hO����|n�1|s>�o��x���7��M��{����������'�Oy�/���zm�/��G��/�{�G��{�3�c�%�r}ڏ��s�=�����_��1��|���S_�W���O&�ϱ���'�E<Sޔ��好�O�^%��_\��5�g����^�/�\��r>�����۵=��?(/�'~m?`|C���l?@yi?���1>#�i�_�O��_,�9��O\���~���j{���ƿ|N}9��g��|����E���E��?8���������w�?��W�����'�������B�Ӿ�����C>����@���;f�C���_;�/�7�����Qm�Ƕ_���W�o��眏�S����>���0<����=�x&�l}ڗ��_ߪ����|O���ƻ�o�Ϙ{�o߭m�9���i�^����33~���������/�����?~�}�o��X3?��u�>�߫=r��~�l�Wk�Oڗ������������//|�1����6~����ܟ�?m=�������A��'�wg�����7�����IQ?���nj��/ڃx�<{��S�?�K~���;ڇ�r=>�|���ў��J{����ڞo|�|J}�9��=���k�{U�g���o�Oyh?�/�[>�ߛ?)?��|��-q=��S_Ƈٓx���7>�}i���?9?�F��-�������������;��s~ڋ� >�/,>�O������������Ɨf/��=�g�Q�x�s�����V_�>\���������}���^��4?s=��rm��{�� ��ն~�>fO�?�������;���s>��O�X�N�q��i�������퇉7���}���/�'��{����2�������k���������?&�����'�x�?��/���p>��:��Z}`��i��������G쿙}��'~i��p=��1}(��_�|��������oj�_����1�S_�o�6�??=������x��m���7X���+�=�������o��|����oն^���~|~wp��#~x���/�=�o�s����Ϗj�����O��2��|C�R_�����Sڋ����Vm�����E��#��x�`=ړ��֞�b���g��Z��;���+�]�������������g�����M��=8��ē�����6~���'���������S^���������|Ny�?�'��#�p~�����K<�/-�h?��������X����O���oXoŏ�=�e��c�g����'����x���~�|����~���Gy�/�G�Q?���?��|e�1{P�x�����ﭞ���'�3�d��hO��1�5��>�_�O��{��xd����<��{���2�C��?�_��i�D�p�wk����_7����O�ԇ�/��,�Y��vm�[�_��O8��|�O��F<s���?��O�9��x��O��E����w8奿oj��:�_�7��"^h�o��'(/�����Ƈ���_}t0����?�'�-?�����[�C>��(?�g�L����o��>����s�G�Ѿ�\��0���|��-^���Olm���j���}d�7�#���7�[���|���f}���y����7���?@�O}_�m�����~'��H?~O�Ѿ�<�d�����7k�����=�}�����iO�O�s��k�߬�yz�����/�>�3|�}��Z�������囑g>2}~^_�������|��w�����|��!_�ߔ��y�����$?��|NRړ�������C�Q����_�=ק�o�6�t�����ל��0��=��O��ּ�?�w��}�������?;X��Y|X�s}����z�ǌ?���1����>��z|��Tm��%>��E����#_Y����O\������'~hO>�|fO�c������|���>���#_�>|����?��^��i��?;x���o���-��9�]�����S?�O��'�G��� ���N���[=Ky�ģ�G��>�'��?�=�a~3�l?�^m�������Ϲ�M���7�������3����V/���j���?���sڋ��=������GZ���~�|��o�g�K��V�_�/�V�������Þ|>����{�G�7����;t��`��g��Ծ�d��|>�;�7�/��>:x>�7��絿�4��rm��p~�����߮�}�#������}��ڟ'>:S�Wk����}�?|?�#���iڇ��Ym�3�M��~O|����s��oj��[a���:�����g}i�G�ޭ��"��C��~m�>���w���O�i��g�R�i?�G��{>'_�^���3���)����8��|)ɗ�?ף���#�+߷x�}�=�E�����^|���>�c�A��?�������[�C}�?9���>�G��O����n���e�N��Nm�ߔ��3�О��3�q>ڟ|a� �e��~7���VoZ}���7�kԇc�3�����������!(���y�{[������?3�P^ڛ�3>-��}�C<s>Ʒ�3�c�9����s�k�������|p���YS>�Oy���9�|�Vm�K�l���o�+ߧ?�O�Ǫm��~i=g�ڗ�0�oj˟��!_��ԗ�x���6����xc�P�C{���o�O�����9�A�)���3>7~4},_�}�o���������+���[}����ϙ�?��y'�]��ߏ��Y�s�=��'������z#�x��1�[s�~Z���Y�Q�|�y���s�w`����zߩ���<��/��<:Xo������~Y_��o}����^��Y>���{���K9?�I���/��]�ߋه�H���'ϊW��pL�[��$�����{��0���|��s=�;�C>��F��_��<�����?�'����߮��w�>e��h3ވ�O��>����oڏ�������P߁�y�K���O��Rm�{Ӈ�3�����Oy���Zm�K���|�˝�_�ը������z��1��\����7�h����<��C{�9�������)/��||N�r����c?��i��D�#>)�e��e��k���W���ByS~��|N{r>~O��{�����}��Ɯ���s�C0�i���V��R�����z��I�,��>��|A}�9N�I���k�����7���σ�����O�'�m�g�>�x�~�7�ۿY������|My�O�����|>�o�8?X�E������k۟�|U��#�S>ڏ����'�a����>�G��g����K���_�~�x���>�EY}My����O�R~���G��?�j����=��>6���^�}�g������}V���}ԙ�(/�S������5ۏ�S^�7�1��y��|���������#��;����?h/�O<��C|����||��~U_���?o�v?����������;�z�G��6~����'�h>������W��
Gx1��ߌ/ڇ뛾��+��_�����S>y��|���O�G>�zw9��ԇ����ߧǟ_�K}i?�'��s}�G�9?�O�߫m�j|Oy�?�/��Q���O<�/�^���Vm����6����3~�<�������<_�ߔ���������㻵��7�����g�%�1<s}�+��Q_����|fo�������ƌ�+�g���?ԏ��������X~%1�P^���C�����x�z��2>�}�?��Mm�S�/�iƇ�����K}�/���g�A{�|�x������ ެ�!Z�C�2y���z�o�O�^6�iO������ߔ��7�1�oVr~�!�#_��6�i?����s}ڛ���������O�[������7VO��ԟ�`����~�S㿗k�O�z�c�/��=Y��}L��a��j�����N�o2�?�1�ð��_@��>����y�_����7ޯ���?�=�����Z�������?��Bm���x��_Ol8����z���nm�p}>��9?�9��w���{2��}�O�O�O|R^�gx6��ԇ��s�G<���'��8x�1�#~؟a�`��������9����|��&�K��}6��f�����=jK���L>�~ߪm}3bc��s}�����|�1�Ϲ��g���\�|N��|��]�ݍ6������È�:����~[����?&�I����Wƿ�O�������(���s��9���7�7�~?�����9&�џԇ�SށU�;ʷ������x�~�_9?��l�,׳|�1��x�|ʱ�=�Ky�=���y�������;�G����b�^�툏_�G�������/����c�~T��~�k��O|�������|S�ϗ�ϙ�D{qL<���g�a<�{�7�IY~b}A{����?��x��\o`c�=�ٗx��|��#�����O˧|��'����?��s��o�ǜ��Z�l����9���7������@��aߏj�m����������ާ<������j�~~�Zm�ӯaߑ�������/�W���ok_o������)�	�#X�0���vs���k���P�_�6�(����g\��6|�x��	�;�������y�jˇ�?�����o�������O��o�v���nk�{&����_�����O���x`|���'�!?�Z����1���ԗ�2���7u_���o�N�����|���|�3�=��O����f�ޮ�y�o�H�������~�+�����&��������~|��������0|�����_���x�sڋ�S��,�������qL~��ԇ�g>�|@��oĿ���g�1�rL{~����f�ك��������/���?ߜ��'��/������l������m>���oX=g�4�c�!މ/�����hڋ�p}���?�u�ڗxH����<'^��y�K��i�g,���k����wk{�k�������)��w9���������"�����~�����`�_Ծ���޿�-ކl��䇵��Y�����Uo���=l����`<��|1�'����Vm����?ß�_x�7����{�`L{��(��ws0��i/�o����{�?o�ק�\`s�����}��Fm�����9��M������'�g�>�O�qL��{��rmχ��O����Զ���M}��><_Q�{p�\/��o�G��o�6_�}ڃc�Gy�����7�����ᛃq=��}��g�O{s=���s�û�+����ěه�o�����>:x��"�������Q���R|������#�����'s�7����iO�?|=�k_<��><�9�#��s>Ӈ|;rvT�>��#~��m���������7�'�'���!��7����{���g��?,�~������|��f���qL��~ć�O�=��|�x��,����_���1�#������B��}G�z��9���zV?�ϩ?��F���ߤ?�������9塿�/��G��?s>���_�g����=�O��ǘ�x���4�=�-�3�a������>���f��5��<��G���X�p�M>�~{���o�o���r�Gd���s�o�˜?��-��~`�xaj��'��}�����3�Q^�O{�?�׶?�nm��q}��>|������盗��_�'���G����}����G��I|r>�G|q=��ex�����|f��j���=Z��2~�?�#_�����1�'>�O�'~�x�~3��W�������>��[�:���qL��{ڗ����?����?��q}��>�����I�_9ǔw��/����ɴ7�_�6��ߴ�e���s�N��=�o�o��z���<�׷�&��ԏ�����;�������w��7��b>��io�3塾��W���(����A��}��/������W���ն�o�����3���������#^:xN�Sڟ����j߿��qy?��ˣ���K������������zVOq}ڇ�0yY/�O�O������^į�GY}k�7�K�h�'�'����on�O�_�����1�Gy���������� ��o�/<�/f{�wg>��������?���棃�)��E��g�����~'�����?�y�,��7��ٞT_����̷���3�>�m�w�Ǉ�X��7k�O�=G���޿;ҟ�����9�W�z����>}�b�n<j�/�񈇙�>�}?u������ߧ����x��菛����'���Ԟ?g�S��<�����?i�C�>�-�q}��c����'��_�o�'��~Oy�>��������z��ڞo��[��T�/��x�V��� �����=�7��s�{��Fў��>�My8f�?1�[�g~��"�ӿ����������{DG���B|S~�Ƨ���K�X~{����K}������$~�>�I�S_�+ԗx�|�'�g|��[�c|B}����ԇ�&��/�G��rL}�^��-��9���|��L��#姽�/ړ�Q?�c������}�[~O��VOR���96>�|ԇ�?�wj��{�׻�m�M{O�����N���K����|K<�~�/��z�_���_�������Y��x��My?����Sx~�����'�����%�B{?���_�?ߩ�~��?�-�P��a���?�{0��?�_c�}�`�=�cp��/7��W��?���)�?��t`y��|����7����:�<�����{�������Q�/x?��}���O�?���)��2_��?_N�k{=~������O�O{Q�����5�o�/��0���?��_�G�߯m?��Myi�Wj۟������k�'ڗ��/h?����W�������?���o�W���y�ʷ���I���c�������G��އ�ퟘ��/��s>������Uړ���X���s���g<�9��甏�s}ڋ�z���w��߬��S���M���O|ҿ�#��s~��M��V/|NqL},?R?����M?��Y��?�1�0{>�-�=�K�$>�/i/��������o>g|�����:���?׷|G}�O/׶�K>�?�ק��ڋ�r}�C�߳��=�ԇ�r=�����;��c��Fy�/��|B�;V/������~�1�����)���;�}����m��~o���໰'׫'2����}���~0~\����b�w��0���������7����́~#���5})/�/�v?�������F���N������o����z��?�/�1�5��.�C��y=ڛ���h/������ϬG�1�w��=�9�ޯm���P��Am��k��a?�������ԏ�?�����}�<�/�K<�^ԟ��||�|��oj�/��->��K�Pڇ����1�w�O(��k|F��X������X�|3^�/�������~p+ϣ��	�%?[����}������\/S_ڇ��1�D�Ҟ����~��ǵ��r�:�o�&�i�ף�������ף?�=���M>������>O����ޗ����ȷ������hx~8�����S�3����=9�a���������F�Tm�|��`}d�3�g�}���7���[����g<�S���S^�=������x7~��M�S�_����������/���������ǐ����߯j�?{��緿��~d�=̏���Ԟ/�������<��}���a�7���5<��G}����>��E�������@_�OR��k>=�G���ɷk_1����ӟ|��o�ψg��X�?:?�v;��b�>�>�}���G��9����k�{�>������|�������|N|Y[~��x�s��K���|N���|��~�?���?�����z���9��矌�G~b��|8�_�g���������9?�7���8�x��/��x�|���Gē��c~�?�=��2��O�sS�����~�k��/����W�����S��ڃ����'�ړ�R��_Lc����ޗ���O��O��>��x#��/���=���1��O�=�K��־ޟ�/������ǵ��/�������3���Y��Oy�_)���|�Ϧ�凴����/�c������Sۯ�~�������Ɵ�#�����=�k����'��P�����i����k�~���\����[�_�~�������_�;�?����?�k��U����������=�7���}�3?��m�����2�y���1�{T����x������{��>���am���׶@�>�����������|o����?r4ߧ��{~O��ԗ�%>�0z�<��������޷��X����������O<Ѿ\��q>�~�������c�ڃ��|��[�ݟP?��.��%��H��G>c}��ֻG�&�Q?�����k�e��ȟ�w��s�K>�� �w��@_�;�a�3>8����/�O���������"��=�M��>ăك�H}l��J��^���}P���������i_�㦶���x%~�w֣#�������:�Gԇω�ǵ�����>�}�>�|�^���ϩ���o�����~��� ~i/�О�ն~�����rm�}1�����Y}K��b�>�"_�{ڟx�����C>����ǵ�����<|����|w>����~������y�����a��?�/�z��s�/k������^m�������g��j{���~Y�x<�w���񼎿��}�y�������wgy��������(��z�Ԗ�(/�!�ho���G���o�_[>|ts��ڞw<�m=2r��|�/ԇ������}x�5�3���ߩ��7_�����ǵ͟������k[�?ԟc�[��S>~���G�g��!�����rL�pLП#���$��/ڃ�Z�O��Q�)�B�q=�|0j��E�S>�G<q}�3�E��/��c~$>)/�sLy����}�[�x#Q�������s}�Gy�/�u������������|B}8���w����}8����s������������m���3>h���������Ѿ|����|�/�����#�ߓP����`����ϔ��0��}�c�x\���7�O�|��f�2~(�����9�%����+-?Z~�lL�����-��\�� >�o���������o�|V�h�jۿ��=?����Q����9d��1����Y�j[������o�y�,������n͌�ٿ�����y�?}��}��>�G���~�7f{��1�'�Xb?��{fy��g���|�z����ko���>��~���~�����/���!)?�����cևs<P��g�3�<���"~�/��G.�l�\��6��'�Ep�ǵ�������?����9���#����������b��}>�}(/�'>)?�3~���'~��-~)�i`y�����7��M���#�ok���T�W���xb�R�4^9����|�����Ә�����O������:��hO�!��y�=�/�!G=:�r}�w[�����9��|��E~��8�#�h�o\�����w��|��'�7��O}���m�9Ї�s��j������C����!��?�������w�����������ɚ3_�s0���`=>�z���(��a�a����`���O����7����{�>�}�Gy������qm����y�:������~#�x����<|1�3���_3?�<�������|�k���?��������<�>��`>���nk��)<�ƌ~Oy���3����7�=/�~R[>f<����^���z��A�9���\��B��/����G���j�����G���/�����?�ߧ�9&��_ȇ��x����o��:�g��3>�o�'������W�O{o�\6�s���y\���ڃ������~o��������w`���S>�u`g޿2>O���#��ߧ|a���?�wڋ�r~�)?��o��C���q~�z����1����b�������K�K{r}��]ާ�����Fq��Ծ��~����/�1�K��9�I|�>5<��S��;S�O�P^�O>�<�k��K���x31��/�����,��;�5�!����C���ǵ~;Z�O�/����{�����=��o3^�~{p��Þ��ٟ�g�Q��?��g����e���%�y=���s��E3�����|��O�s~�3�o�W3?��$(/�e�P~���1���m��}7�;X�������ev �����������ͯ���}�_��|5�?��n����{s=f�F{Y<�}��)��{�=�n�2b�����A����1�׸`r�'�E����7f>0�^�z��2�#�)���A��<|�.��-�0�����]_���C{Q��{\��zƋ���0<�>������O�~��߫��1�����s�����'s>�CƷ՗�'��$�����o�G�Q��:ο�˻��O�}�G0�3>�>�s�������k�/���a��s���ڞ��~�~�'��R�����Ig�Fl����4���E����<��{��������҇������7���oj���~s���6>~����|<��)�G{����G��,��ǌ��־���͛�6�ߟ������U����)ޟ����Ym�������������)/��s�?be��?�壽�_~O{>�}��_�7��Ӟ��|D}�g�O<P_���w����)/���ԇ�`|�9�Dy�����|A�����x"�>ף�>�m�����-�#��|�x�����ק�L>�c`�_D��O�7���큾�o��O��7����0^�?���sL����F|���_�����*�q���x�=��>��}z��'?�����V��\��E})���%���`Ԣ�<�?)�Ջ����},^)�mm�?V�0>Ɵ??X����V��9��L�i?��l�߇:�/�����_��I{�\��&_X���k�����=�oڗ�������31>������_�ȷ\��E{�����|�笇��>�۹^����k[���f�猏ao���<�x����t0�Mm���z#����p���ϼ���'���|����}�Gy�|�q���O7�xp�3�?���2�a�����|���Bm����������y���#~�|@|R���q}�7����5��~	��G��<����s���ç�|�7����O#�>c?a^���>�/�'�_ڛ����ߧ����=����#~���>��1�:�f�R��e��ŌǑ��o>��mm��#>ȏ�7�G�O����\?3_���W��~ԟ��\��f��o���b��w�xp+������h_ڋ���'k>k~��|����r3�?�?8�����ӿ|��ܿ�|B|0^�g�c���4f�e��o������ޯ����x#ߌ?���9��a��}�w<�Oڛ��|���J<p�x����xb<1��'�Q����^�'��xb|~R���Q�����ߏާ?�_�o�k�˾Z���-��=��<o�}5������K����ԇ��~�����~�����������ܧ��[�G�y0?�|K���My���ynk��'>:s}�G�G����7��׳���G���<��/��Q�ff֟��7��3�s��o��#�Ҿ��f��<\��q>�o`���yL���O�h_�������y~����ϩ����������O��G|q>�����e���O��Ͼ�o�/<o������>�{����s~�t{�>�C�h�7|?�+�?�I����f/���nk��\���0��F,��`>�-_[�Y������:�c�о���߿Ҿ����{�#��?������'������^ǜ��o�����#�O}韏k�?�����c���1�A~4��ԗ�ў����i/���(���^p���߮��N�ӟ��x�?ު�}C���w�?�g�~Z=B��oy�n��Ζ�=y��'�����k^��`>���j�o�7�������zo^�O`o�?���g��1��;�Q>�O�F��ϋ���~��ٟ�����������~?������/���3�����חk{�N�~�}��>�������ߩ������G���[���Y����7�g��U��)\��}^��5�����q}ڋ�E>e���?��B�F~��>=x�x����sl�O{�R��[���on�c�J�>��~����_��$��F>c���?�/�����m>�m=L����/��?��O�-��ڏ������?���(/�r[���1��2����[>�=��c>��|����O��E�hO{�� ��>'?�=����������|����|�������W����V�0������_�_����?���k����G��G��{�կ��������_M���>���ؘ�����7O����Ϡ��9�����t�w�O���6�o^?Xo��Ճ�~n�񈽹��}~Z[����������������g�%�g��
��?���i�3x�������9���_���|��Y�m�3�C���3�\���_ڛ�P^���?��~�������[���+�������_������C��ߴ?�����o�#���x���?���f���6bk�_)/�7�/z����/�C��9&^��K��^ԇߓ�8�ԗx�����6>�|ԇ�#�O�磼����x�˷��8��Y��c�o��I{�������5ۏ�B���A��^���'�?|N{�R^ڇ�d=B�3�hO�����9_��ŧ��1�g��o�>��V��������8P���_����x_y�����G�	�����|>�?�����f���{���]?��������Ǳ����������|��菱_�{��>#����N����޷`��}����u�>�}(ߧ>��x?fΗ�f~���ԗx�<��A�R?�;���{f��em���S����>�ާ|����g}�O��&������ެ�}�g���O���%�'��Ǽ/5�K}?�m}�Nmϻ��ԇ��3��+��<�O����M���o\���>��=�>��c�O{S?��G|���>�Oy)�N����>����?����8�O�p~>��3��'��۵�����c�;�Qs���x1<���ߨ=��C�_jo�g�a����??��������z��Ay�\����������|�O}9�|��\;��8���K�"��>�~ԇ�����O�����m��3燑/��i��|�~�o3�������d��}���÷�_���ې�o�񗵏�e���+�O��9׿U[<q�����r������j˟����_?��~�������7������H�nj���?G������S����+���?�m�;�a���k��a|r>��7�?ק}�ǵ��c������9�e�G����7�G~�}�Y��k{�� �8?�#�߬�y9��|߫�}������G<3�9�3�X��)�9�|5������ԗ���ɚ��K�����'�8?��}F��}w�/��H�i/>��̇���/\��\:�e�o�>��M�y�m�����ړx��q�7�S~�O�R?����{G|M>���?��������3�K{R�����a�����)�B���g��o���7�����1�K{R_�ϟ�w�=	������<����o����s��I��c}t����߁��i<��7�_�y�<���۵�G߯��a�C��>��߈����=����um�7�G����|1��i����Q��|?�����?�-?����'�Ɵ?L�Q�p?��l����������׈י�(���q�_S��o?<xN�hO���A{R[o�s�qm��/k���}��+���9�'^�����{����e����[�~\�c�O�Ƨ����{��>�M��|�3��c�}�ڟ�o��1�����9&�iO�3�g�"��~�W��=�����2<s=��Ok�~^��E<����E|�/��Sڋ�By����9�������������m�����9?�������#^��\�x�z����ğ�\��%��_ն_7���=���?�㐟�����#?����}�/�}�Yޟ¾�����z�3���4�3���Q����߇����D�(?���� ���:X�����!���Ay�f|��������#y�����9�������;��o��?s��|@��o��;��́=�|�˜_F�����棑~|0?�?������%�(?����}��ǵ=Ϣ�)�>b}���/�'������>���$^hO�7�M{���W��K=��}�r}��������O���x\�j֟��=��O�qLy�_(ψ���|6�0��Gn��Q��+Ot�O��|Hy�>���io��3����:�����-(?�Iy�?ڟ�"�/ק����+�G{r}�kc��7�G���G�S��?������3����w�������b>�z��Ϩ����~�,�_����qm����3�q������>|�k�o�����N�����~�,��k�a��ό/�����[X?�Gyמ?x�f^��͟#^�{�Y�������_������c�퇵��v���9�i��>?����>�cx!^��������7�?�d�_߰�?�7�7������\OҾ��ᜯF,��Rړ��^����s=ڋ���i��f��|�+Ǐk���>��+���4���I����3�)�#������w�������O>"h�������u�����'0ߐ�����>f�r}��|��h_~O{�?�V��iL<Q_ړx�zԟc�G����ϴ�}O��o�c�O�#�2>X/0�iOڇ����oG����l�i~O���|�x'޸����������ڇ��X����j�����c������#�� �~_�x}��g{��|v�|�_�/g���y~0������ �|���7��b�p�������̗\����������ڟ����s���y��1�����;ާ����p=>�>\o���ԇ�x�9���ӟ����oj�{���,�n�'^�ߩm=����mm�L|Q��y~8ۏ�0�hڋ��>���3����؟��jm���j�ߋ�>��oj��)/�Cy�w��E�o߯���>�?����fU�/m�Ɵ��ƌo��_�+���џ�ק8?���L~���o���G<��Ư�������x�|��c����?ԏ�������m�C|�z��>	_2�Oڏ�|���_�> �/9&�R����\���}�ړϩψ�Ək�?��1�s�m��֞?o���{���y�ǰ��o\���e��=3>����;�L<��������<r��?޿�}��j^��~��|�v��׾ޘ��=�o���~R�����E�}�����|�x�U��<�ioڏ�s��j��i||0&�?��n�=
�W����~��/�����|�����~��п��Ծ��=�7ǜ�|A�����o�~��Zl�g�+�J~����xe�_�~�/�w`�i����{������0}>�m=D�r}���������/��/k����)?�!�����������'_�O)?�G~!_p=�K����'�C�0ߑ���ٗ�w��|^7����ޫ�}��k�߻�=���My8�W��7��oj����1>��7��@��������N>%�8?�?����Q>~O~�����Mc���?���H����#��}�����a��ÿ3_yf|yXOr5��g��g���Nm��ǵߟ�x����~i����ǰ�́�|>�m�o��c؛��~|>�?�˯j���>�,�j���|#�����0��_W[~�g�o�o�ϫf}������?b��-s<���)�y��{����='�ޔ����Oy9�}>�m�3ꁙ��O����}�>�<���Bm�m�;����`}�7����Q�r>ڟ�Q_����k_g~Ny)�#_��L?�K>�|_�6>>��J�ҟĻ��m��G|K{0��O��x��~R������'��򓿉?ڟ��|Ư���9�;���������!�iӏ�'�R�Ok{�F�v��@>���h?�����������>��=������O)?���q���B�y������/����nm�������s)?�'�hO�c��O������H{Z>�����}��|C������)�#����W��}��_�>������_A~�7�5���>��̷ܯ���ߧ}�]�|��9����f���W���{��Fl�~�,?��1�EyhO�����s=:���8�k֟����}���?������^����iL�R_�O}������"�K�>�m�j䣛iL|Ҿ�/���h~O}�O�3��qm�}3���u�o���p�k��"�F~���9?���?|���}�?i�Q����q���C��v^��������'2߇�y�/�K}��OҾ�G�3����}���������'�(?�C��=��W��/�������WƗ��+�A�8�G���R_�����D�P~�������+���s>�G>��7�?��<��1<3��9�g���������W������̗���>�X��/����|���i������v�����Ǉ���hk�������S�Զ�����~�|ߊ�<���������3����o����k|>�1���}����>�~i擁�W�|�*��{�Y�G{�������ר-~q��=�2��������7�������1��a|1>�����~�������y>�K~�?i/��'���W���~)�3����c��ާ=�����?��%���_6����+������'�����x�;�(�ӿ��������7ß��O�2��=�G��o�����S��޷��xi����~�'��G�;ڋ|����]��x�����O0ߌ������8��/���7�ߗ��xd=:�g�r��^x���<�~��o|?��������{�9���x�2��5�=�g��v�����ňO�Wُ���O����f�>�����6�ߦ���3~���"�/�z��c�1��\��?�������?��z|N{������;���P?��'^�/�����?��́�|n�g�qL�3�^��y�`��qp����|�_��W��o�s��۵���6������v�z#����x����g�y��Ŝ/�oԏ�B>�s��;���@y�g�G{0~h�����c���)/�I��O���������������z������y�l�N>���7��!�a��:������^�?�'������^����#�V��@>�G�ؚ�����/����;���=�7�=�����o�����\f�����a���o��9~�C�������������k�_��k�'ϻg��~|N}F���<�;�7�O�����x��)߈ϙ��8��)/�������;�{hޟ�}��{ڏ��;�s�a�9��y���}�z�+��}��?��������/2�?��|??��r�G�p{�>�~���/�'��l�w������Ә|3����yߟ���x����>������1h/��G��9����{��������������x"�i�C}�?��3�1����؟��7����>�c<��?�I�S��g|q=ڟ|D���?��~��?�0�߭�q��4yh/ڟ����O����^ԏ��1���(�՗���0~�w�|���|�w���֞�g{����7��O!�W���!��Ym���?�m�����ῷk���|��S����~ߌ߿��h�O�W����}�y=ڃ�r~~O�h���M�����G���qs�=��������������c�����������#��~��_�v�B}�ӓ���3�Ϲ�x\��Y��'��w����G�b���]�~���x?���,�F�Ҟ����(/׿����O}8��?����1}�/������������s}��c��������=�������cޏ�ף=����}���j{ߏ� �����@^�����x�?-^�/���~ԏ�B�0����8��k��=(/�G���ߣ��_����h�o�K���8����C�����������1�{��i��1�3����/X?��[�����>os}F}�X��|3���sL}��f�Qߑ{�xx���G����[��J}��x�?8�8�}������Cy���j�o#|v�=����OG��z��Ef�?�׶^����`ޟd=��W�����3�i��-R����x���/�O�ho�{�����?����'����߈%ޯ������8~���_�}������?�C{�����{�s>�~�o�^�9����ԇ듏�'������?�ƌ��/��?�����`�r}��Iy�o�g�='?1ި�E�~U�x���_�/�E�О�w���i�����Yy��5�������o����F���Oa�����?~_��������|ß7����H��?����)�K}��=������#�.�~~��5���9�;�3��j{>D�R�ǵ��|��ڟ����>#���`�d<O#g>�=i��i��]���Әx"��_����/�?�O|p}�?�奃�V�<���G���烏�z��@���6�C�䣙��'�`�����/���%~��Q�����v��Em�����i�Q���o`q�7�����_ڟ�����?|=�Ǧ�ԟ����{�'��f<���o�Ɨ�_/��s}�+�?�_�G> �rLp}���6��g�1���G���Cy,Y�����g����Um�-�O�<�/�?�������/�OF>��������~�<߈Wޗ����=�2���p�a���c�؏�������~����������D})?�7{Ӿ�3�^���}��v�>�x$���!�~[�z�v��~b����y?0�cη�ۈ7����I�~������#�C�S��}�Oc�������k�������x��(�'�����ԏ�E�~Z��x�zs=9꿹>�/�����������Y���B�~U�����Sڏ��}�㶶�M/�?�O�����O|��/�K��g���ڞ���W����i�wk{_��e|Q^�G���|���9�#__�3���gӘ�FsL�������w[�x 0(�6�<׫�G��o�8X������} �8��؏����_׾�����9~}����~3��;�����m<Q߯j�������x�����È��|�ߓ��x����?����������3���8�+���|qs /ǜ��ڞ?�����^������;��<_�������n���^����?�~�G��W���s�|E�������{������������x���,���{��x����<������ڟ�O�[���{������?>��>{����|#������> �>ԟ|Ny�w��|��g�xp�M�Q�����������_��ǉ7�;���)?�E��zv�Z|�P�i�w�����G����-����;�o������s7�'��l��?ߩm������,��g�/����#>g�����a=3�\����Ϲ���g~N�G���5��������x>:X���o�?r��R�x����-?�x��?�ی?�a������?��:�:��Ey�g���Z�>|�Q������~��?#?��D{�>\���O�o����\o��\�P����끾���Dynk{~�����s����G�c����q>�'�K{��ԏ���#����k�_���[��x�?F~���x�f~N�>��}w����}U��p�����|A{R�Q����m�F{_�Ϸj�O�<�?�����/�1_0?P_�3�A�b�}Y���{���1=�m�x&_�[��G����߃�����ɟ��'ߍG=��.�h/�!��� p=�k��֟�������z���nk[�%��������������s}�_ao�?�4�ǈ�/�g����a˹�����ѳ}F����'�gy������#>�������<����O�o�k��k��o�����n����>�����>��y���������B|�����3^F<�������������{���Oīً���)��G�p>�����1�!����A�r��s>%ߍ��OӘ�O��<��|��{"3�i��s?�����>���5��s�F�߯���L�kԓs}g��}iO>g|l��4&���+k�K�9�IyG~��5ڃc��K|�zf��^|��g��8�������������3�]�����/�������8�5�W� ��|4�1�{��\6�`��e~���/�a�?<��os��O��������g�=ϣ�_���C��7��������j������i/�O|��5�'�����#�f~X�����~�ϴ?�%���3�s��;�����Qg��{}��>�9�N�_ԟx�����|��i?�7��Ӄ�W����c�:������� ^?�m?���s�k����*Ϗ��1�C�/�K���}��#ߎ�:�7ڃ����o����3�g��o����z�ԇ�������9b{��ҿ�o\�����z����(�હ�0�����?��Am�O�_�������__��\��R�G���6�~�{�|�����~m���j���כ����+�9���`�;�7��\o�����1���9Xo�����=~�{����X�x���ۓ������c�{m���<������~����F���Y�~\���W�+�)��3��\�>��f����m�|ߕ�����A{Q�k��</�}�9�|#��3�G���x{��>�g��k�'s��~����=ڇߏ|4�/�O�Ҿ�����k��O{����|�����k��}+�e<ߴ�e|<������;���>����ϧ1�q�3�י�K��~�v������������4&���������?��O����?�/�M�����	���������Ϩϻ�?zvO����r;��}���f�F��|>������~�����w���G���<|��k?}�g��\�����l�����g|r}~O����������o��c�i�'��1�3�鯁Uޏ��O�Q~�?��+������Cm�u��\_��x<�ǟ�e�����x���.�ܷ�Ok[oԏ��x�`L{����=��鿯j������|�Fm��#ڃ�~�����_���x�䕃��'ԟ�3�����?�����o��C�i�_�������������?=X���u��|N|q~>g<�o�>��s�?��sڛ�1���T��ǌo��|K��[��j�gܟ���g����6�����_��3��x��Ək������9��|=�����֋��o�������0�9���@^��ڟO�`<�w�~���n��;����2�cp�Oڛ�����^:����|�����/#>x_n�����8�|ԇω�?��Ӄ���m�a���7ڏ|0be�K�7�y�o#������/�����~�?��+��W��+���~P�~*�%���/�M{S���h�7�Ӝ/��QO��h�~��Ə|N������=�7>�?/�'��Ip�Q���;�����i<ꑹ�X���z����ӨG�����ϴ�C|��O��Oڟ�d|��'�7b�˃�ǟ�ہ�\�����/j�{¿������D?;x����O�;�g�Ӝ_F���c�K�/����}���i��u���>����2����Y���/�|�_j���xx��K{>����-~?���|���>��7�`����槽h_ڟ�����y_j�ǈ�<\4��(��7�>��w�������'����O��o�?�������s=����	�O��({0���\Ք�G������@�RIMB�� �0E3HChi-����!�"����z�c;�����*��{�ڢW�׋��{�*y�w:'��<��W����o����O��nվ?4?����I{��2^���<���#�SƷ�=��O�[�?�������/�Z-_I��'������U{~+�}><�o��$>'~�x�zޏ|����J>7����o�ϊ�?�|�B?��<����4���l�E:����K��h�E��O�;��w�g���_���x��ώ</�������z�cr��G�_�jx�5�;�=ϫ:���;ď�y�3ǟ�����S?���7|c����y���gƧ�|���N|�2^R�Q������~�����N{�����9��״W·|������i�ϵ�O��?x����%?e=k��=���<��~d<�����s#����oR韩���C�G�7�I�I�+����%�%ަޯ��p�C�#��|`��oR�����i�|^�I��|���G����"�F�����x�|��������r�=.�=s=��ß��5�W��B��2���ߺtD���W�;��O��١��c�#���'�T[��vW��\��c�o�W~����/�K�7�G<��W维?�?72_�)�A��{mz[���s�'ǟ�OK9�mo���x������ī�'�)��F>4��~s�Ŀ� _(�k5�b�L}��?��|����'������K���?�y���|6��~�>Ē빜O�|;+����������x&_%K��秾��]�������'_�����u�����������S��������C��|x������?�}33�R_9������}ܣ�~[�O�#��������=���?1������k}1׹O��s���<����+ߏ�����_9l�|)������?̟������?��y���/����̏�k����,O����5|���ý�_�y��>���_�G�+���|�~\���������9������_��6߁�=d���Y��S���s��=����W����O�?�7_-_]�����9�T��E�o�;��σK�?�{��^����gd���O�L|N��|��oW��s<i/���9�'���~���z��#�Z�x�^��5:�����6r��ؿ櫍�C5�?���s=��O�_�o|��7�������Wm�>�Z|ǟs?��	���'�Οx����S9��/�7+|s>�o��������2x��e��ě�=��j�~Y��}�Vo��������9?��?���������N_<���>?�!Ǜ������x���Ձj�Y�#�w����_P�?�O����%���S�����|�2_�x���~ƹ�r�/�������j�+�����?���5�Oi����=�/o·?�_�e�?���C}�|}>{�L}��ˌ�oy=��~��/�v���j�g�[��ܿl<xZ���߇?y����ߣ�|�����籾V���Ģ���x��?����,o�#�%�������r>Ğ����9���Ϲ�E<�އk�>	�<��~�C�?�������x�y���F��Vm<�=�}��!��߶W�����]��ӿr�y�A�G������I����W�?�'��|�J�a<^�a?#�i�?����I9���͟S����O��%վ_9�O>0>��3��5�m�7�=���x��i߼����'������>��ė�K�wt��Gb�ɒ��·�k��C~?����]o�?��e>�ϧ>?��"ǟ�����H}������_�/�g������'r�����􇌧�~�g�/?�r�s^g,Gþ���j�������ԧ���1]�!>f�������'�p�-�sx~�A�K|��|����>���7����������W˟�k���۶W��t<��s<�垑��+��oN2xm<I}���wi�����g��|+���wc[�������c�����������|I��Mr~i��W>�|��2/�_���Ӭ/gG�㇯N�</푟O�Y�a�<����1����Uk#�K{�������O�j�]��|����������^��9�ė�~>������'����j�����%^��s��?�/1/9�-�C��3ǟ�H}%>ݣڿ�����`݃Fdr�^��B����xB؃�9^����b~ģ��"�W[��'����_V��X���^#�s|9���*����ި�ݣ�^�����?�����[>���?�~�����'s~�s0>�S_�<���;��K�����\���^^�?�O�o��K���G��?��H����9�?���g�#�ޘޯ���Q9_�g��_9��j�3����g����j9���C��%�������_?�����x�\��7=�y���\OO�L|�w�?oR����'�i��w�i��_���]���W�o�9��o�?�x��M�H����x2�r|�)����?�ܟ�σw����j��*��E�濧܁�����~:�н��\��K�_�Q��ŵ�s�����]����^XC<q<�/������/�����o^�ޚ����^s�)�}�5�G|��+����G���xJ��xҟ�/�#5��;�������s��o��ͷ��O�_^������Ɨ�O�k~>������i��_~?�=��z��"�-?�/�s��o��������&�A>�~�?���?��'�t����B�/���?��������}?-�~g%?������>��|�N#��������~s����_����1?{A�3���O��>�B�/������#����v����|r�ē��o~?�O�f=�����������o��ll~y=�s�ֿ��KF�~��M�g�ZN9Ǔ��g��?���|�G�#��P���&_����yS�/����O�K����}�^O<�?����9�ī�ϴ�/�5�����x����-��|,�;�C}��!���8?�/���p}�׹��������s���?�e>Or��������p��)a�C5�{���Ǆ}�_�G�������S?y�|����;��8�0����l��k���4��>����B��S���D�?;�ݧ��:���N�����<?��'��\O9����z��xw�j�����O���)�$���R��{~��V?)�O���c$�W?�W�#�g���E��~^�K�'�����r�7���5��{G�Q�?����r�����_�O~?�g���o����f<���������~^OK{��3H}��%'>�Wk������������o�/��><H9ǿ���r�S~��[��|���~y����������W����g���M緧�=�<��x���|�T��/���'�O������j��u��x�O�$>�yV�/�������z����ώω�9���`��i�'e�)���!��8~R?���g�'��
������|ߐ�>�C��ӟR�^����?�������G�Ç����\��3���i�|�b������o^����|x�|��O}�0r��^��_�j�'��/��%[���R߉y=�x����H|KM�'�9_�������ć�_�O�;�����r~>��9_>�|���~G��~�_����|��/�{����_��v�-|����?K���S~����7���#~���+���{���j��#k�?��g�_~����~Գ�ϳ�쮖�����o�'�C��x��r|�[�K�W�3�3"�߆d� ��Y?M�|�x������~�gT9���O�9߂o�y~��x��]ɗ},s ��������=���<�_0�g���S_�5|�����_�|t~�x���/�\m��K����y��|�祬�+j��\�O�M����w�'������zi��H�/�s�j�#�����9��/�3^�5绌�GT�wO}>3���/x����7����7����Io�W�������G�|>�)�1y�*�I����R�|w��Y��~���G~~{������9����_�_�����#�����)؟f�ldۿ�s��F����$���<��~�/�>9��GH�\/���Ǵw�/��������䳽#����xҿ22~��i��G��|�ML�N��ϧ6��W��	����u�����̿�^���w�c�/�>�|��K<L������r|��i���|\��X����3��~�5����^����Cnw�,���|��Y�m��5�W�D_r?��A<��Q��s�;RC<7��1�����)�/�������.#���c�#�Pm����_�����7�?��3x�z+Ǔ�����o��xK�9�r>9���?*��IN��Z����Ϲ�l{��Ɵ��'�g����o�S��y��xrY��x�O~>����'?>`�~�?x�O��5|����I�H9���O�ߨ��s���Y��7��|wqD^��߿u�H��|3s��_�������_�k�'���j��$>�=��QC�g{<"�~����<�|����z���뉡�)ϧf��B|}���Ї�;��[�!~e=����	���W��_������b�=#�ߨ����e���X�;���_2�<����0���>�����W�~����>������1�C<��j�x�h���O��Y�/i/������3�#�_�����������5\ϴ?������D���򩌟K�}_"x��+������K>�|��I}��?"��s|�G��ײzhD?i��oڏ��z(ǟ���3�s�ċ���5|_�����1>�Ws�х��^���k�������Or}��{V�������_o�kV2����<���s���M}������2>���Oy>x��#�� ��O����v��k�?��#�'^������x7_ _?�G����{���c���^ù�#��R-�~r�O�6����7�����Y�#�#�|g���{%�/��^��'�C�繒3���y������>�9�?��g�3����~���g��3>s<i��N�����I�x=v�����/ٿ2������9���{揌��_��+j�>&����_9��/���=�{���ul��oO<?������7���]�^���3?���c����o?�����q<oy��#����y>Xth����|=����s������y^ޏ�0��/�L<'>�����F>����ħ�?ǟ���_S�9�Wl�{.�L���+$������7��ݪ�C��&�A,?Nr���j�Wm���ת����ϜX�l������S�Z�����Z��<�i{e|����Z|M���=Q��iy���O{�����T�����/�0�������j�/e<��3>Ӿ�?i��k�>�{���|x�����x�0_N�%�/�`;�����H��������O��~���x|Y��'���6�]����4�{Um��~�����}��������Mk#��K�xu���?s#�'�/�ϼd���[�>/e�?����p�}#�ze���1����?�~���<|���c�M}�U�7�S�~������\�-T�/�>��秿f<�~�7]�����/�3^6��;9_����������gJ��?�x�O���W�G~??����z��~4��\t�祽�^o�Y��Ï������������6��C</ϳ��5</��/�Ϗ�.W{�	���|�}�s��^:~�N��9�}^��~�j�zz�~�|s4��M}����C��:�ar����'����Q���"���O������ُ�pD���^����g���T�{�����?m�yG��������)�x�R��d�o�>�y��xQ�zV��|��{��wO�v�>��}���}���S_���G�ý|�����Vm|��3����#�!�̯s��9燜O�/?��I}%����m����W�gC2��|�)5|?���aծ�<����=�V�������p?L�������J����_����Gy>�П��n���z�?�3���xc<�����x���R���r��<�����e�4�oT��`ϼ�;W���^��w;����'J�^:r�����<N>x����~s���$���k$��p���^�I~b��(Ǔ�_f%�W]�f��wy�������oy=��K�N����{F���F�����w�7Ǔ����=���R�o�K�?�_���|�V���o]l���H�o�o�7�'�73�o��<��g����43r��j���؝�ZO�񿲆`_����9?�/������Ò��c�q��1�\�����た��./���o�N��z��s��+j����w�'�+�d�yp����x��g�g���-�E�8����}��k���t����ϡ�ǰ=Rp�9��K�#����x��6�^\-�������M�'痟OJ{�>����G��/����C������d<Яx����+�7r>�}��|%�3����K���/��/������~9������_�/����xA? ��_6���~o���{��o��6��ί��x��1߼~(�sY��U�����O���z���w��<k��rɬd�����S~i؇���E�ߗ��^[�?��k�9��U?�E�/���������#���̓G���M���y��)����r��x5����ϴw�xc�"��<��}�����y�}��xE~��t��s?t����/�>򕒉��zh�~i��缞���I}���ο�WT�ǗW�5|V�1�'^�x��<_�xL� ��Ϥ}�?�6>O��O���χ߉9��j�'�k��^�[�o�/�(��K��O�7��K��/���*����_��?�?�k�����}�~�<��#�J���������g��2?}f����o�x[~T�;������=�;_��p����b� o_��+$?Ə�V�>��%���?X�z/�G|�~���yp�?ǃ�|�d���\��狶t�-�����N�J�����#�|�|2Ǜ�ϲ�<+9�~����I��o2�<�=�?y>��d�o�ﳿ�x�z>�%5���罪�|������jX�X������[�z��7�s����'~%����N������{O�a<��\����k}�|R�Ү�祽�o���|Zm��r~'�9�s>y��j����@?&�;�~A��$^���_���|��6��s���{�</����O{���W�������׫i?�/���ȩ��/�}�9����9W��x?�jx|ψL�5ާ?����Ӟ���ٓ�q��e��"���̧�;^���^oۨ����0^��cb<����kj�~Y�,u�����v�~>?�?:�W�K�?��I~F���a�+���\�����s}��K}�|��{�</�ω�g���W��9�����x��ܟ���������_�����������<Ƌ���#�Z����H� ��JNK}e���·iߍ�,�'��{F���x}m�8?��������|��N��������O���O}g<?/���9~ȗ�/�ܰ_~~af���C۽�m�վ��h̏�:�r<Ŀ�?�eS���%������~�d�i�������?���+�r>J��}�|>e�۞�������N�@����N}�w�_�+���!=��U��o�%�]�7��q���r>��oΟ��ۈ|��������,1����כ�����������K}f|�>3�s��ó|>�����j���:�ƈ�4^��Q:�����s�&���/<�������|���Y�7�5����[����ϔ3����_ӟ����m��~�����Z�~��r=��$o������Z�W�������y�Y�G�>����5쏺�xz���Ǟ_2�<j����y��z$��������όg��5/�^՞�L}�_�G��i���r�N}���W�?׫�$������c�7�jj�~�|�Ɵ�����s��#�3�zu�W���Ӿ���j�#�-��H�H���UO�����?���`E����C��\��Ǽ��|�$�^ �^�ד�������=���۱}7B_/���M�|>������e$7B����A�}�I_m_�7�*�G���r>|f�7Ǔ�Uߧvو�m]o�_�����=ǟ��&�̎�3�~?s����Oʩ����x�|���������W���^ī��H����s����Ӧ�ҿ���Gƛ�O<T��Cʩ��?�%��I�xK}�?���ί9��ׇV���g������1>��x�~/�}�:�w}���ﮪ��?���˴����uy����j�9�x����k�~I�]��J<��6�o����[�n�����ۧ�ת�w9~��ղ����x�g�s��x��L���d�O�C^�Ύ�_�J2��������2�b�O�Q_��Ǖ��/9�����9�W���i?�9�y~i_�����o�<��E��o���~�k���"��-��?���j���W�i/���0������}���SN�����ĖNl�ԧ�����p�zN<�j��u1>������/��Wא\"�y�/�cnd|�S��]G���������j�����#�ڟ�>��x����/���������s�ܗ�\'�w�<?�O~q�}�����������#r�+�������]����<?l9����C#�O������\�|���R��?���#������y/�_��Ob{^r����#���,r�������o��e��������������x~�W�g��O��~O�
�5<����xf�����@oY2{����	�P��'���B�����p�|�a�|^��)a��9��{װ��&�w�J�����3'�d�K}�o�Oio����!_�>[�߿��|��'�WU��įׯ���M��7��	Ώ��WR?y��V臸��'������ �^?�����W�o�C�/��~�^���U��4>���z7��������z������q��s�7�;���O�IN��_���ŋkx�|��5<a��)��U������ˍ�_��}�M��`��x4����G����/���xZ�|c���������xh������=�<���9=^�E��s�ǃ��J^�6?����ZOI}���ȯ�G����k�%r�������y��/x�|��|h���Y���=R_9��Gr啒�w盜_�;�+����[���x$W8���,T���;�</���4���͗3�ҟ��w�U��ӟ�y�}�o�����_�����Kkx���ﮎ\���=�g�|����G���w�����'��;�y������ߋC_�����>�h��5|��{�Z_��7K���<���|��G>��K9�>��S_���Xt��?��G���gݶe���5���N�x�+y����'��?��!>��i��W�#�o�H�����S9���x�|���� ���4�"�ޥ�;<�?~�22�����p���7W�� 6j��Wį��Z�M���k�ۏ�s|)?�Z��m�׾���9��'�O���Vm}_w�4�����+~��xe}���=_ě�{������a�'�K�8>��w�<��.~�����&�:>�/�c������������;~��|���}�\�O}l���'�C���y>�y����?�O}�<r?�5��|�{���9���,|��2��^-��/�L�0��W�o�x�v4^���_޼���������'��?f�:����^Y�L,������ۚ�L�1>���`������ă��S�^9ޔ�%��������䣾߱�'��m�ka[&_�s������/�����xw<��ٯ��r��c�_�?�_�����w���|�|,y���r��Ƒ�����������G�lz�d�5�3|������j�;�����6�5��|��m�x9'�|�O}�ƿ�f�����wy^��z������ċ|^����3~>9�1�5G����1ƿ&��t<�o��+�>y��5ܿ`>75? �r�V֣�W���L������?���۷�����	��?��=�����ώW�vd�ħ��h�W`�|\�|$�G����d�;\-��茶r~��\���k^-�x7��o�w��'4r=������>��G�]�w~|2�LY��~��wK��:V-d<������i��|���%���S��a�W���ħ|~�S�G�'�)�߇��I�J��|�y�����_�g���s~i���.�`k��W��E�|�x&>���߈��������s��i��_r���'�]<�y��x�>��~�~x�|�x����#��i�%�g�J������ƃ������S?ė�ıj׳�����l<H}���>"�ߎ��/�����[��K��O���v���q��5��_�ĳ�xw��W�y��o�?X��e�Po_�Vm�y������<{ľ���j<9�����~���_�u^r�ӳk����?�_��^��9bqnD�y����j�#��)���/�W�{�w_��yj߷b}�8�\m���L,=v��ă�~�:����oΏ�7��G���q���b�o��^V�~�������7���j�|t��Yy�b�!~�?9^��|*�s�j�K�=�k�<��?�n~��}X��g��d��xL|��M�<3^��6����7���>c�>�?����;�w���`�O��_�/O��o~����_;_�������#2㛓������|�k�����a��M|���Ӊ��?�����es����t~~h��b�����e�Z�����G� ���ޑ����:�N~o�_U����ot���%�����/�i��g%?�Z|���>!~�Or|�E��_�w�Z� �r�ٽF�G�d>~�^��~�?9����֫���O��<0 ��<y�'�9�Anu�"�oR��՞G<�����ěă�W�A�~��/��K�������f�a�+��?����a�/��#�ǿ�6�}����+kx>��t�:�N�;���C�������������}����{9��j�m�|</��~��_�/�>s����d��� ^��+Ə7T��ɏ��O�|������S�_�;�3Sm�.�'�����)���������ͱj�wH�o���</e}���#�����_�X�ԑ��}R>_|����ّ����ȏ�i����}�����淧��_�{߇i�A�y~��H~��l�p���~��_�����1��^�]����~��k���}��ϩ��2��/�������r���ǿf%���'z3o��+ǃ?�?�x�_�ob��d�b����?ҟ���������I�������x��L��O�g��G�_��b������_�>�]��r���%�p�4��|�����������<��z&���j�u��[�_�7���;�xS�y?r��e�|��������?���s�%ߗq��������o�~��bD_������5<_������'�g��5>|��&���j��B��`y��s~���<_����o�c�Z~�?9�xRO�6�/�k���.�����;��ǜ�Ҿ���6>�E���3?8R-ۨ��r���)���'���9��O�O�/�^�������������9W<���G�����������w�k��~O�;��d�n#ׯ
{~E����ϋc~�{�1���\��׈���|���F�i|'�\�⯳aO��Z�����/9��x�1~��S�9^��[��o>W2�������K�A~�#�x����S__[-�>�Y�?�_��`�˚Oܻڿu�Z>��#�:ߥ�o��8����$��S������ۨ���%�G��]Z�����_h�����پ���d�c^2��|�/:��9�7U�)�g�+���{E���2^���7�o���x������G��,�*�)�_e�x��$>�_���g��O��x���ǹj�>���#r�?��<t��i���+��M�����s��|8������u�"��_���D�/�+��?����������S-���������|��1������k$����j��C��w�j�� �d<A�����ч����w�x�����c���j��}��u���_��|��=�_�9���e��3�e��I#�#��$S�-H�oؿ���#2���;��q�ݖ�Υ��k�~D�;�����7�tϑ��}��\_��8��������R9^z��VۏH��?�����|��x�����E��=�?��k���|(���O��ʘϱj�~1+>;�1�-V˯ȯ޿�<`D�2�{y������4߻���pב��|П�EΟ�����k�yy�c~D���|Rr=���?r�G��y~��7�</�K<��7�m��4���s������?�x��r|�g��e��N~r|�|���۞�����'��?�~�͟s�+�~���<�����7{G�o�e<>'����0��ԑϣ�\�����Xߏ��l�O>???�e���yj�s�Z{��_9��>��Z��ο9��/�"�G��t����襁��j����}��܈�R_G��[���<p>�����W��s~�����<�n{��?�w�#�O{�~����:?��S����?�7���|������������;��z�|2�G���������e����9_�y�����'s���9�������+�>���'�SX��*�k�П�~j>>���]_O�|��J���T���x�[��s<���nT�?��ߟu|�?���_>�|�9V��K؞W�p�����~����$_ۿ���#����|��� �4� v�o9���|xd�L��O�/�Q�:��|�/�i��k��a�H�d<^Sm�>�1����[���>;2��x��`������N�����o�O�ϝ/ӿ�~���s���'��#����._���_ϳ��G����a���k&\o��������ӕ5|?d������#�㿯��z����'�5�W����������?��z9������/�/�Q��"??��\O���mGFƟ����}R�k�>7��v���O�~��7�_�\2���=�y�����s#�H��>��s�'���x�51~l��x���&�I��.��^W���K�����c�W���7�Wÿ7���F�w�|��j��P��:�c�{C��n����?���3p>�����y��Α��?y���#�s~)�U�/�������?�O��;�/�_|�|8Ǘ�O��>�[��_/����6�������i������3�����^�"��e|����i�;�E�����r���R̍��k�~���_�}u�{|��Ǟj�5�����v��7��w��ē�)�j�xn������x<�����ﻌ\?\�~Y�b����{Fd�����o�L<��o��T�z=�����Fd�;�/��mTk�|~ڟ�c~�������K�A��W�g�����zϛx<�_`S����|��'>���#�{�G�[��|��K{��ӟS?i����=�]?I���=���s��x�� �t�yO��EЯ��_}�~����|��+F�c5�?��aO������:��"��y����|���u~��Z<Ɵ:rp�^Q-�_̯��'���C#�M���Z<���r����{�#Ǜ��^L����s���u����=�ǿW�<�\�~b���j����'������7hw��c5<�j�9Zm&�>�~m盌��j��R���~���L������;�j<oV����k��̿�/�/���	��������?����m�/��x w>o�����#2�l|%~rH�����}Gd������������j����L>t��{Ɠ��'�~oS���W����'W{����[��������7K&_�������o�=���|?�>��6�q�����K&���WԐ�Y�O�����?߇i>o^��v�y!���G=�&�5�'�xc|��9������ל/��׳����.����Y��W��'<u>���/���/�O��������S�ީ/�3���2r=����񤾈_��������S���P���?�������J~w�L�Ï��i_���+�+�����ٖ7j�_��;�c���^Z���ٿX�s<�o���O�y�d��� ?4`�ϫþ���G�����/�3��?�����
����Я���5���������\���_��s|9���^-������r�}����>���S��v�������+��������>��x��j��9���$�w|�������/�W�����r·����ܯ�������w�7�����罦���="��j���w����u6.����+�G�������7���W�������'�����s<����G���02��x�=3�z|��z���ړ�q>+�>�����u���盪����t<��s�y?��|�s<��Z<L�{\�����j����Y���c���;�����F���R�8?���F����c���W�+����U5�d>���緯��8�yu�U�!���#��|~����c�筡��=�����Ǒj�ӵj���������E��R?�j��ӫ���'��q>I}�=��ƿ�-�l��T럩_������/�E�R?��\���s~��s��8*<3��t<��9~�E2���%��7��x��^[-�ω��?����9>6jx~wo�g6�o���x��Y�s����o���?�|�=G���m��|s��9����~4��C�!�)�2��s?���q}���_���F����{F�������s�����#G������u�����Α��o0��_�ĳ��.�o�:��*��x}���>����?�߱��|������{��v��-w`�}�_�$������'�������}��\���]Um�K}��;!<5ަ=��u�~ɖ���Ư�O���z��#s�i?�+���\�C����ķ���ě�C�;���ڨ�����%?�Z>��"�����pE��+B?�ϋY_Z��kX�~Bד����������/������/�=��?�r��U�/�A�Wq<���z�����k�2������>k���9_�����_W�?��gK&^�g��3�>9���i�k������'直w��|�������{><3�J�H{�=�W_�{��e�����wNr�C�'��>I~���O0?����=�C<;~��<o���<��~�5���`�`=k�������x�f~E����ա�;W�~�?���'ǃ=�?��Ms��|��~w��������O�y����~�zn����2�>���j��r����>�G���=�}���n��-�_����_~�mDď�)���������ҹ����gd��#�O��'��\;�o�g���8���a���X���������-1����5�o`�%_O^����3�y�������a��?�?��{���7���x�ZU��:��F�o�p�����ş�?i/�����µ�����ȏƏ�'���L�j�7x���֫�W���߼�Z|M��?ۉ�������/���o��������M���o_�K���#2k��O����Z�'�q����ȿ��kj�~ʹ��9�9��}�����o��k��z��E>{�_�W9�|�?�/��x��]���o�����~����5����\OJ�c�N����_9�c���k�������ư����������/������ճG��u5|�������Z�w�'��f��HK^.��5\?��֫�{A�O~�C2���$�k<�2?2���?_s�i?����g�oy^����*�E�;~�UO9�����/��S&���:�K�����2��x�#�FƗ�M� �r}�������~�;�G��!՞O�;�P�W�p����~���3$S����'��?����_����7r=e��� ^:߼;�.����f�3�s=r�����{������x����?��/���&�wM2�;+��|�����q磹����Oƣ���×V{��x0�?���s���������%?\6r�xr��//r�i�)�+��R_���<���8�u��D���k#�=�������L����x��͎���5\r|}M��Z��o��7�y|�#r>���?�ח���xv�"?���}�$Wm�l�G������~�|O�|�d���x��9�?O�/�cڛ|�|H,�NT�Ծ>���3�[����]ڇxp���y;���xV��O��l~��;^���?X�W2���"� �7�����~�m<��W�9�,�?�_����~�d�aN2�ea}�|�X����JΗx���:���|���s����s?p�O�7��9_|�%#��#�O����|�wU{ބ�m�zb���o����O�z��>e�!����0�ϱj�|K>�������o|K}����?��;F����̗^�yW�>E��\^-�������C�|�xw�#����`��#�'����%�t~?����N}��_�(�ߟ����?�G�9�/�3?�����u���8�������?����[����7��kj�~�q����L>6��~������~��K�[~��j��X��:s�i?���/������~k��Q�c�'����a��5|��������7nT���>_�G?��_��kkx���#�|�d��������~`���v������#��'���#��|:��/S?���x0'�x�?�o����g�>����)��?o�_��|B~p��������������5�1�ٰ����1�w��V��wb�{���a�g�$^8r��a���Ǘ�)����������w�'�$��^<���_��x������x ��?_Z��V�go��O���?�j�O���G�O<9>Y�4�K{���Q�y������_��O����̯�>|��2�Χ��!|�|,�9�{;^��<�`�^���Ҙ?��z�M5\��^�y:�C�ho�/�ۜ//�6>^��;��w�/�7��k�~���r~���=�uT2���x��q����?��kÞy����9�>s�y?�����s�~i?|��k�?ǫœ��6�������?��r� _q����k�Uڏ|yב�y?���������q?�zlV2x�x�&��1���#�;�=V-��x��ī������6�o}��ѧ��3�-�M}j<C��_���	�q<~�ֿ�Oڋ�0?�\��ޚ����a�����K^_��|m�3�C>�������|�r���A�������#�%�������7���=���|���|uHr�?xn� ��l��G�tx._�_�o�����o���s�x7~�g�?��q?�7�]���c<}?�3�a��;C?�|�oy����{$��_�d�b�G��<�??2����j���x�?e���L=�����Y����������\䩒ɯy���#ϻ��z'�����c��$_�>^-'�>`���j��`���+k����^�}�y�s�ó�2�u|��{�|�x����_�����<������z��J�co�o�c�%S{���+�_B��Z�F��?�?�7�����?�^9��~��<j��o�_b{�|�k��`�J}��[m}t�6�����^�7���o����2�%�~>,������9�g�!~�1"��Y-A��$��<�<����55ܯ����!?͍|�C[��s� ��:?�}��|�����N~��|xˆ���=�7�c~��S������ͬdbﭒӟ�Ϻ��޻�-�W�%��y^���/��2���c�u����������G��8^�_�0���7�(�z�d����}������s�O��9��_�ģ�M���C�xk�����
{�x��=x�x�o/R���O��ˬ�̷��=#ߧ�h~^8���Wķ�)�����j�M�?�������qE��7���?��o����?ȟ�OC?��E~��)�x�~�������/��������~)�<q�t]���ٟ��v}{}��{[���װ~��П��*ƻ�/����D�y��5���5�c�ͯ�?��觸ߜ�*�^����2?�|�1�S��ܱ��W�؋��oD>V-?go�ɑ��o��5��0^�8"�?�=�������H��Y��z�/��9�&�����/Ƴ�	����_ѯ��r<a�\������K��-a���>9�����/�S�?�ç�����X��o���6�|}����ߨ�Ӟ���oڇ|����o�ϳ?�=��Fd�ߞ����Kc>����ޘ?����W��X���!�g�"����\���v�^2xi�=V-���O�7�G�hV2�+�A��r�!>�'��%__ÿo���7��i�+�?>n�:��G��$����y�p��K�?e�#�����G�+���j���W�_��O8�6B�o���F�����z��Y�i�Z{;ޙ������p��͏����x�^��f��ߍ��o���R��W����L`����K]������^�/����5^����9~��a����m�����9���������C�?�E��x������#�������#���xe���2ާ���r>�?�o<z]�g<����|����|b��v{ml[�8�ȏٯ�~��яl��xw~�_?����A����S���5�"<i�������^8��U����o|��������g���!^<�<���r~N���k��Gi/�b~��O���2�wO9ߍj�>������z����O}:?}C�#�/�~>��5�{�6O��4+�Xp��]�?�{�d��F�}��6��7·WT�9����j�|b~�?���O����j�t]�����+���5��:^�O������K��5#~��ī�$���q?te���7��R��c�_��`��;��|��{��/����+�7��|��?���'������O_�/�܏|g�$>O��^Z��~��j��¾�O����y������w�o���$����������z�x��Ϗ�~� �x6�����߬���M�F�S/؟N��啕>#~��×�|>�=\/��O�?'����g�/���5�d}���6����<��S��|��������z�����f|'��I&��Oģ��x4�}᷏�?s��-���>^C|����~����=sw�_6���'�Z��/���kX�-��>e� �p��%���kħ�ӛj����o���=aO�����?�~���>f~��R?���|h�������|p��}�0���s�����WIN�#�^���U��C�����'����׋��Ώ���E>��b���?a?�O���rU����ׇ�ȏG%���g�������������w�˞���	:���� �Ӽ~؟������	6�;���G>�Q-������/��i�[]�ώ���<�a^8�o��|9�O�2>�G+#���z<V�j�臷�ݖ��]��O�x����ć��!_0r�g�>���pW�VF�O<υ�o��}
��z��?���#վ�~������?k|��ïFdb��3��R9��+��%�����>/����Z�$�/�לo�>��I_�k��v�H{�������/�7�2~2����G�r}�����G$�y�y~��9^��O�x�+�I~5�ݨ�_��G��7���߰���s}�ck���{~����h~�����W�U�#����������Z�9_����g�������,���;�k���c�/��]G�G�?|���-�;�pϑ糾�~	x�W�#�l�����Ɵ/Xr��>���gT{>~g'^�_'jx>��#ߺ~����'t}���_Y�~���~��Z�~9?��s����99>�$ï�/R�ħ����xa~v������Y����|�G>?z���H��G�����z���������ғ�}��l�g,�����+��gt�~%���U����������������7�~s=��r�E캾�_]_�ƛ5|��x�7r?�Y�OO����|M��E<oR�y����_���u������|��m��Gm�r���uak������:?}K̗���=f��p7��P?8~�'����}�ωj�}.�܏x3>��ُ�}�k�𱵑�ேF�E~5L}�O/�L�����?�=����<?��r�E#�O���s~���d�����-�||p����K���+���� ���W�gڟ����Пxp</�':�>O@��{�yĻ�	�0?@�����������3��z���|H-�c�~��L|���/����oi��S���������l��K��k�^��ҿw��~W�����wD?�k�����c������#�'~��'j��������v���a?b����νG�7�}ѷ�������_��o{|����!u�������G�~��pc��s��K��=����7lO�����q}@}��	���~a��_S��E�cď�#���x<V��m�+�m�p��~>xi<������'�Ż�W�`w�׌�%싯�?C���z�����z���5#��W���y^��a������7��x~8�|S�9��'������_PO�yL�[�������w|��6$�G����7��~̏��Ϲ�I�����w��[je��D��o���O�6~�.��z��ߎgλ��g}172�j��u�)��`�/��������5����<�����r���6~�_�/��|�&|N�|���?�x1ޤ~���O��϶|E�������M�������=���ě�5�Ѭd����;ި���=&���L|f}��=���Ɨ�~�Wo���{�y
�k�<5I�Q��/�?G$�W�G�����9��>\�����?�1'�d�x������+��K������)���O=d|�p��l~@|�?�����sb��c|7T�W��gI&��o��3^�+���6�V�/���d�3�|_B�7�Q?/�_�?�xs>����{�W�o���7���!�O~���7XR2�k<�����W�?��xy>}���O���9^��x���I&�IƟ�w��c��l���~�ׅ�X0��'���j�)��#�����1��g�|!�I�?���|����<�����j�+x�����m5|ߑ��<~��i�c��#������G~��u���@>q<��r�N���x����xh~�������Ϸ�}���o俹���K����7ߺ��|�~1r��N��I&�=rnv�d��#�?�#���d�_.�~Η���#�Ş��t���o�u�w�����;�߉j�!������������>�����p�&?�V۟D���ׅ>^�������ģ�7xn|������^2x��y�+�r>�oͅ=̟���R��ϑ������!���j�k���ww}s]\o]��_)�4������;f��Z��'�e���=O2�����'x�xG_�߫k����o��/�o�W�������W�;|��%�	�{����U���r>)�/�����L=���/x����W��*��2~?�?��{>�d���W|�e�W�t�-��O���|��w׃��������T�__���_����7ǃ�$����'�/7����X�w�zƹ�G}b|�1"c?�)�m��x��	�<�_�?�e��\����O��o�L~�~��E�+���K���·i����x���~��l�kw>I}�?Ƌ.^���L=i���������yk��>����|�����S[:ؖ"�}�Z|�?��.l�>�I�7\}U����{������r�O��_[����J&�?���wK�?[���w�O�O�}���?�K�r>!�y=��[:7���{�k���3���x}���|a|N}���_��;���=��%��|��>�/�S?���;�}�kV2��|����z���~�?��#��6r7�e�&�{�d|�`�O���G�o׷ϩ��O��1��o�����%�G��~����|o|8Q����O�W�߄xu�%?�K�^s|�/r�Ro�����Oi�|���OU�w�Y���X_���I���B|��\/��������������������?����?�����	�K��|�Ώ����Hm��'�G������/�+�g����}s�������ڃ�����t���j��0^��O�Xm=L>I~�x'��?����?���ǵa��~�~�G���j�Q^��?�J�K����'~$S/��$�WF����Z���_�%߮oOV�����:��a#�K}��P�~%�����V���%{y�'�o�x_���??R���z>��v���Z鹞�����x'����\_�F�����X�L}��
��|��|)�����O��Ò�_������9�ħ�'����NW�^�� ���I ך��^-�j�g[��Z���Z~�o�/���������I~A��X��4��¥J2�8����Gk�^��Q��D�x?p �K�����v�]���^�#�5�8��������;�'��6���u�i_|��K|�U-�����w�G�&~"�3/�y��c~ԣ������T�W�xd/��\�|�ڰ��z2�s�Z|I��j���u��5^��?�#�m���?���w.�����k|��z���m��7r�������>����9�ĳ��/����xM}����:^��|j�!�:���瓌����� >�$�����/׳���s�����7��2�6�o�W��'��$��?�׸��=�?b���B���t��H���|��㛗_s=�Θ?��r�����?�}~�xD��������ߎ�q]2��|tc���9�S'��������ˉj�	s�៹_��$~�/i�_�{;��k���S�x��z���}�3�r��������m���|�����ѷ��t}�~2�'���&���Kվ/�t~�O��G��WW�9�_�6��W�������~���+��̎�?��K�1_����g�7����5<�`}�]vK&޳?���탾\߾�Z���K&�簷��ٿЗ��u?<�y,�����y�55|���u]ϣ/�|??��H}�_�/����՞G��M�~.��6>o�?�'��p#�����/HO�$�r�I{�u���u��7��_�2>�o��1�C|���_,��C_����|{,���d���m����<����/���џ�#��j���kx^l~D?9^���@�p��>{����/�h��ny>��Q#�O�\[��	�>i_���v{m���x���Tm��8����G>��j����J���~��O�[�C�˷�p���~��_��������Ϻ^���'X��Hb������i��ߜ�r��B�)�a���&������W��ݖOU�oė�w����I��џ�x��}��~w�'����7���`=��#�9��<r�7��~����9^������g���[���?���W�yN2���:�}������[�/�w�Z|a�ޯ7��Ϝ�药K��8���<�b��/�>"�m�o�`_�3�����I���?�4��߼�yվ���x#�ͷ^Z�~Pj�	xl���j�9���*���F|�O�~���<6�����r��Ϳ�7H޹����}]�|q����o���e�k�W�_#���~��9��F���ׇ�'��9_�u~D'�����	�:,|�����3�$��&�7��﫫]?"sүK�1���܏�vِ�:����7z�����~.�o��_���ڟ�W�?�'�ke<@��*���|w��ް/���0�;�%�G�O�hD�?fG������:�m�?_NV�W������h�듩������
;>�߽#ϣ_���������^����O��C�c/�?��3��6^?������>�}�ɚd�_x�/�s����#��������~����/��� o��������O\��ϏW��ă��6�l����<]����=��_�Wr���v�KΗ��|�t��������a~����C��E�#���#�s=������4��1���=[ۗ�����|�/s~7�=s���|3�sM�x}������O�1>��\����x�8��x���7�{�d����鿘?�����_��t}H<���?b>�����7���0��_�?�����D9�W����Z��4�����c��W���j�m�;�ji�/������!>�|C�_�g���J���aO�7|�񏿻�Ŀ����9�����xɟ���O������>:���_�������r�����F>���O��n��ɗ�����a_�=/������\'?��>���?����x�~M�G�K�_\����#���<��L���^�G>��j���5���;�C���^�_���2J��9��O�O����#1^��z�|d<�?�7�;��¾����:��#�>���_�~��a�#������Z�����j��g�|:�w�����ɏ������|��x����}�>�k����>?p��/�?����|��8U����o�RO�O�/�\2�c|�^�7x�|H�a��b�;^m|�U��5|_��<2��_0�~8����/��z�a�{R���~����kx���x��;�A=`��������w�m{[���y=�O��B2��|C�w>��Z~�?:?�v���̗?U�?a�K�+�_�����aO�����e����|����d����x�������������/���Z��ӈW�+���Ώx1����ۜ?|�������1����������j��&u����g����OZ����	�j��{��O���G�O?��c�������j�����<���[�t?~�罍���t�-Z���ߪ�^�r����u>a=���a���������^?R�������џ�*ǟ�������'�b|��$�������������T��O�������?&?:�?.�{�>���������d��+$_Wm�F�ƻ¾y=�O~��9�O���"�wc����g>Rÿ�����J������/�?�qC2��?>���z��I<��w��6f���{C?��;%�^�ގ�(�����j�p���%����>�����^�����������_���B��?���=r?�o^���������~��/����m�?�_Ώ������/�|"�C?��K�0�E��������7�O�?=^������g��bo�K�m|�8��׳�����9��Ւ��wKK�K�������|M<���?��ێ�o�?����-H&���}燴?�yx�y��7���d��>�G2�m��M���C��T��n����<�����G|�I������j���=�Z��f��3$�@��x=U�~������K�>(�����ɗ���g�|&�c~�z���D���1���E�3���ާ�������x����g�������|�E��`>��C^o"�:���6_}(���%�������j�%���-x�k��o�/��x'��'r����;��x����~�σ�η�����xB���~�k���ʑ�O������[��{���ƞ�7r���z�d���y���7�/�%/�O@-���{�`~���>B�22��?x�x$��6�<������|����۟�W�O�)���T�'�7�K����J��_����׆~��ۏ�|�_�'|����1������|��j��ǽ#�C���/�?�����}F���~D2���}�/�u�K���W�#~��|G/��!Ǔ�=Y-�������T��7U����j�;���u�o����1��ŏ��1^�������<a#��;r?��7x��&�{�ό�?��/�����|�ߙ�?�k������)|{N2���;�b�9Um��}�;�v��]a_��~����߼"�����O�xOV�����j����̉j�%e���|k������+|��������O��L��O5"�?���?$z������?�'����F���;�O?��sS�x~�Yop<}y��a�&����Ԣ^��~����~t�Z<�D���jx�����lH�_r�'���������c��;b~���.\��3�_ٟ���i�"�|#�h�zJ�ޛ���o�ß]O�O���?K�q����!\�]�����|��4�oۿ��d���1~�+��+������d�7��}�{s��Y�o�G�������������Ŀ������K#�Gy^�����~���Q�i� ~�OXO0��߮~4��=o���V�ߣ�v�B�or>�Ǐ����������_����|��������x��?��x8]-^���׉m����Y?��_�|��{����A߹�d~C.��d�����?x��џ�����z0���t��xi��������SG��F��lo���{c���x3ހ��H��|d~���O����^��Ṿg|o���c1~�:�o��?�����_��G%�g��	�7���Y�s���f�����s}?���~������#��'���H����'�O�Cs���^��^5���/�Y��������WJ>�۸?����Tm<�R���;~����&�~���B���[����^���#l�~%��x/�����_w�<���Sm}~��|�+�1���e���<3�����{L����h��߭�NU�R_�7�/ÿ�g�ǂ��Q�mH��A2�n>H~q>��j��������'kx�ʟ�L��A���X�<|��H��������I��~��G���������wJ����b�g|η��d����0^�i���+�kK�!�1^�w�?�Y��s����|���Ƨ��v?L���#�þ�$��\���8��o��$��؞Tm}���烷����̍�������S���X��ǫ�^�����|�����������\��{���~(���a�����a��?��߿V2���O��c���*��?���>��r>8Qm}O�p�������/��#��n>�|��c|�'�V�~J�4?"�>�O�g�����E?Q����zX��p��|���Z<a��^#�ǿ�G�O���c��䛫�?�5�������1_>U-^������ɇ�O�^�����z#�(�k��l��_�����1^���vc��|4�@��s�����B?�ħ������������w����G����GNW��o��߆��o�X؛|�~L��%[����~����ǉ/�����ߤ��)�e�I������_�_`�1���yɬW����;����?��o޻�!�@�b������x���3��o/��Z�o0����]Wm����%�Pm=޹>����?��>��>y��u��xWp����'�ں����s����\g����?8���G/�A��z����/�]�Ǟ�/��|w<c|���|u�����xu[�����5����GC_������o_U�����}��3Ǘ�a�ƃ_�Ћ�f�������Kf�^�ĳ�����Q�?w�xs�@��>��7"���K��Z<ŷ̟�W8~R���Ç]�/�^��q?������O������~�����Qm�����k�w�i|��/�n�F2���|y����w�C���O�'�w��~��k������t����#�B�k����X���[������}��y>��x�����쏧?�����;_c��g�ŧ?��~��n��}�b����
��o��c�_���a��~����F��c5�{�'�����w?���1��^��?�`�������O >/�>|#�����{�3�mM2x�z����o����7/��z��_{����y�����x�+�C���_����l���_�g�k�/����۟�_����%s����;����s���Fd�k<8U����_����]`?����>���k�zM2x��
�i���w��d��5?S���D|�_�-��L�v�d��x��+�t���������[����e��p��Ƙ�j��?f��??�w�g֞�ς8�����������g|g>��O��ȍ��Vm|�h�^��+|몑��B�|q=@>q<�~N�}�~���9������w�}�������}�/Ƌ?8�����k��ퟁ������{�o0%��?�"��9~�����$ï��@����5�[��#������g�~�W�_��O�����6���Q�~-�+��$�?��S����]?��;����v���<����S5��8�������u����	����Z�����:�w��τ}�Tm}�}�?$~�������}�F>O}m�����G�x�z��j�&���+�K���g<A_o�L>��P���̗ȇk���ܯ����S�����?�i�#����[�]� ޝ>������h~w=E�b�A��O�J�_��ֿ�2��q#2�������ϿI���M�bD&_������z��������+���u���j�O���?���#����ޚ�������o|����q�����_��o��[k��f��Kf}hM2���?���z×�܏�s� �} �o>E�6���������?����oH��?�����j���۟�p?{�|c�������7�C�]->��(��������/����z���?I�����K����_ă��d��r� ���`ϯK&�����7�#�?���>]m�6�����߅�~,�ߧ�`�E���WΗ�����8/<3���b� ~���~+�w[��A��d��x��1ޟ��1~�#����9�<l�x�^��>��|pm����j���w=����s������x|��z��v�O��9����!^\/��6�G��s��C����K��\2��M���gn���w�M�8�П9$�|��	�4�2���_?����7�����G�W��?W��(��.�~�������}T�����/O�����?Q��{9���fG��{��OW�/n�6�S���d�m�?�p=���>�����=C�}͟�w�[�����o�����o���q]��%�1���8�d��wb��ߚ��-���>���j�E��ח������	|����ծg��o���NU�?���x���R&��$��c��}�0_�������Գ�g�m������Z����g{?-�c��?|���k��!��!��1#2����y^���?.>D2��I���x`�">ͯ��'�\��x|����/�d�o�OYOx����'����/��|>��!����'���R���*�68���\�P����kj�ǧ��[2\��F|��_����y���ѧ���?�{����M�����Sy|7V�߼5��w���Z`�Η����L��_����W��i'���n��d����/�x�z�m��GC����g���q��#�O�>����_�? ]��k#2�#�'�p~ ^��x?�gC���U�?�~�u���ɿY������~�s~�V�_'��;��~���h����j���V�|�����/�g��OV���G׿�Ï��\�P?j��]m0a>�a/�������|y���&�<%�;����-1^��������/�����d���A�o��`�ؖ�����#�#^�ģ�|t��G��[�������?Þ����u�G��6��z�<7��S?�G|�_B�{L�w}�ٟї���'���g��ې��?�'�W 6��a�:_�?y��|�\i����z��x�}��w��o�}�{�i��x����8���I�.�u�|���X�~����x��9&��	��'���Ư����W�����������&�uk��D��?r�����!���}�w�~�xd��Oѿ�x3>}����xI?����o�c���O�������'�o뒯�֟ѧ��x�����s�_�K�'=6���~yA�_��`/��g�ޗ�q��*��Gs}�� ��O��^_��"?����~�o�=з��v~Ŀ���������/����+>"���Ò��5��x`=T��ǧ��RO�����
���d�C}���</d<O�C��$�_�?/�����ѷ��D��W+�um��r|���m��C�8n��o�Z����$(�O��>����e���7�n���|̇�R�g�;r�|��?\�}2�Cn�����5���>��a#���'�?�l~G<��C�3����d���@L_��b��a{�^?�k���x���󭒉w��OW��ċ�{���I�����oė���������P�o�<r~ğ�W�Sx����%�_�_u<͏�GF�o�ĳ�����_��?����'�<r?���N�W������σ}�&�x2~O��ģ���5���o���؞����|�x��/�p=�s�|���ʯp����="Ï�^L>����/�	���ο�����^�}�Ǟ��t�Z~�y?X���}�?�5ߦ6r=����'�'��x��?��?X��ů�?ѯ�e������W��su���jx���@,��~�~�k���_�����?8�?Ɠ���z��s<~�>���s���|�Ò�o�K��2���vD���p~_��Y�w}��j�W��߭��?�� �|���c|���?������#���f|C?�'�e~����|[��N<�~)�sc�����?����'��O:~OW�ϩלr~Ļ�:�@�7w� ��_~�_��yR|��J��xb����_���d�_�S���z�����/�v?@~��~2����w�������a�����?�b<�Oٟ��_��3?9Um�*�����'������:^�W�����}�����r=B<:>��F���|��|��c�����w������x��|[��7c~�]���m#�g>�_�!ο�����j�q~?��'�={����o�7�<���B����xJ�g����A����#�/����?��?z�=��|�=�����8>OW˧�'�˿
����r�[G�������7~�^�0r�۫����_�x��7�����¾��}��|8A/oz���������ǭ���/�=���a���%����!����_�3�s<�G���w���P��y?�K��'�����ܟ�����ϝ�������������=�?2__��'k3�m��n:/1q������m�W�|k�������e���9�������^��
�����b~�)�;���A�cz�{8ߑ����7�o7W[�g�;�������wI�\���	������[���η����Y����n]�Wm�$^���o�6��WI��������������js�Ƈ�|�{��֚߂�'��j�R��ߚ��/ڟNU�~M�/�����&���/��٨����u���^/���-��l<O��9��w�~�����������B�p<�x������H�/;_�����j��1���� ^��}�Z�g=�����ۿ~�0��WO��_��!�_����v�Y��S���0[漞������~���������T|��W{B��{_���k���~|�|��O���G���~~�ʏ����C�l<&?�?��&�%���~���y�5����d��-���W����o������/�z��:��|3�?�/��������?���m�~n���j��`>yk��}[������y~�#��5�������|s�'���>_U���q�Z�>�'���W�������������~5�+|�x������[����9]�L5�f��W����ɷ�w��~����c��[�w�U[���'����/�}z��=�����~����������Q���c|��e��O])��~&���N>2����_�GF>O�w|���{����%�o�~p{���t��?�t=��1?�k�c������#퇛 ��>O<�K��c<�~v<�Rm��ϕ��z��k�o�$/�/�J|d�Z��e�������ض?�ħ&�����3Ƴ�W����������?���m5|�����$�e�ې��(>����׬�{>�w�'���C���O���1_���^�}�ϱ����NU����,�C}zL����8>�G�1���#�w�Z<�r?���z�����?�q������'��]�t�t�x��O��	}�A2��x�{5�?a~>{?��~'���O;ʟ}<��H|��:�������|^r���o_�?�5#�����9��S?���ꬮO���_o����	|>.���|��j�9��o_������@?���U�o��f�����W������9����pk�W���k�������������Wˇѷ���51?�o��j�[o��?����OU˗�$�s���1߿i������W�?��7�~&����3�/���/߲��L���$�T��t�#~��G��
���L��<�i~D��|�|���/C��k�+lc<&~��z|r�pk5x>������J&��?�C��~�w����������]��S�|s��q� ��??�/�����O����|xDƾ�W|oo�_�����?�}��#�]��|u���6��W��{��M��Sޏ�?Y/u���L�>�g�O�Gr��o���~�[�~ğ�%���K��I�?�? ��z�fd���O�?�K?l����\o6>ѯt��z���|�d�h]��>����łd���+0�gɇ�s���'��������c|��x��p���>�����}��Y����;�ɿ^��5��'ޝ��^? ^���������^�_��L�E��&��;���:�}r��J�?��o��N~7^���Q�~�r�����[�����z~�xa.��u�5�}S����������'����+�y�Q>o��y��m�|[��j�7��O��냻G��qL2����o��?���s�N}�|��I�5�q�{���7K��u�d���s�~0�G�����л�z*�a����ă����ֿ������@x߯o�����A�w��}?'�|������־���3�/����[���j<?|��g[{��w=���c|ί_��?�������Ϯ����c>�'�����__%��Κd���]o�[��OD|{�l���0�M�������{<�',0 �]?WJ�l�������&��d���1�Y��Z8����~�d���J���~[���}����ߘ��7����?�|�~H��o�ۏ���b~��J�/:��?��|n��S?	O��e��~6�ǝ V��{��>��Ӓ��;�b<�h���7$��̿�g��������k�ݿ_�z�����m�7��xI�Q|��p���`����������|��U#�����c���Z�gb�^�?����x�~D_��Џ㙱����gׇ�s��o�������:�����������_�~���b���#~]���֞}�������A��Ǐ�mǺ���п���y���^2������{x?��~���V}��7�o��4���_���;���ۏ��,������ȇ�'�[�~�}��1���+����|�q}���}a?��>y}|�n����E���ˮ/�G�N��s�y���į���x9!������$w�����ě�k������?n���u�C��~R���Я9���ٚ�������:���c�����C���Q����_���=^�������e������7��z������>?�����;�}�Q>���x�.�ߢ�q}D}������B2�����O�����7�+X�S�<�Z����Z�������\���¿t����}#2���>��iĒ�C������B�T��׏�'`�.}�|����C�߯?�I���Ob<������?ێ��J����嗎|<��d�o׻�ܯ�>t}�t��j׷�w���y���b�����}�����/�>�1�go��=1�/����=��\_�u��>�����!>�߅��??�Z2� ���)��{H����J����'&[}L0w�k�W�tn�?��S�8���C�S��􇒩w]/��篴��`.�����1����Ƕ/�W��?�<��p�4��K���z���\��\�z��Wa�_<��/8��n�=�Q��ǣ�忷������_�S�)�_�����2�����3�ۿn��ǧ�|+��<�t$�g�#��#��Jr��'ܯ�O��5�/�v����v�?w���#�o��^e�����9ɫ�~z���������񓯌���|忇�Y/R���/Zo�����y�[�~H��R=��E�'���ʜ�� ���r{����B2����s�t����]�/6�y��|��ҟ�~%����=�����������~��알��b<�v������m<�������|`���ڿ��j����o�!�?6?z|��;?�=�?���s_������j�˥aO�����V�{>�~.�j������������B.�~@�����1��xG?�W������y�����������w�����t]��m������"���|���@����Ϻ�x���~Xܿ�G=��������|���ǟ[������������}�_�q?��j���=�;ƣ�����y�����/�:�������=�y
��|��v�_������p�L?��ڿj������b_����t�<u?<s�:���۟���~:�z���z�������[����b|ϼ���Jf-kN���Z��>a��_�6ѯ�Bo�5]_�v�|�~������?�Џ9������+�c<'�'���t�7�u�_��z����Sm�z�{$����z��J2��x%�d�l�����\��	]G7��|.��Q}��_	��|��O���G��1^���{��~��zx��v|���h�3�;���Ws<�{����������4��|B��1�'X�ؐ��>�σM�@�zV��� ��z����'�'ُ��_��ǳ����}j�U��>/��j�����Ŀ��x�d���S��ޯ�$��O�����'�|����?ƃ�m��\��w�sz����}l�|w�(���}iY��1��7G�>�H�sL�w�?����RC>�z�xt��}幟�����wy�����|����1^�'}��ܰO2�a���R߻�I�p�^�����g���>�����a]�o�L|x?�a�É�j��O��^�_~��Oo���K����]��T���7����a��}{<�~�K��M�h�{��[�?�ꧏ/�Gr�i]'7�0����0�F��k��j�����s���gn��x��Y￮���s�w���ٲ�����y��u����/�������X�U��x��a��֘��+��E����}��Q�m�G�{��{�G�3�=���:�sR׿8�������[>k�]�9���7���w�������I��/!���ޛ�Q�{�+�����c�>���)|����3�����u��3?���?&�O��<|����/�����6��>��W�M~L2���7zU�����_ޯE�����'�T���ѷ��ޜdb�|bG�.`��w]/�wkL��l�#�g_����(׿���$������z?���I��e�>��/�op���z���Z{��`>�j��2��/{?�šO���xc>�%�}{��|q���;�@_��w�����=�������zO���c�/&~���ڷ�K�������}}����j�W��^_b�����T���a�wн�~�~|�x���gn_'��>��m^2�g��5�������Yz�?$���̏����@�������h����^������yX����9-���xI/�/b����ϻ�[囉�j�;�|����!,��򅭾��k~E~1�i��Ǟ�!��֯z<���~��ӂU�o1_���ߖ���ý���v<�^����oѷχ��}^�:���t�5��V�����sU�������5|��9_m��v����O�?�4�06�_<K��ޞƣW������'��ӛ�����$�[��+����%y!������/������>���O��%������~�?��=�_����p�W�/�����Ʈ�w����?�_���戞wk�{k_������:����w�=޸?6mH&߉o�����.�L-���l������1��y�?^��Gɍ^�'�_6}!��O2xh�^s|P{�?v?�·����}B?�b�c������>������ǽ��?]��3�2�r�;�5�;/��e#���x�~w�3a��'�k��ƛ{��^��߼����۪]��]-�!?��"�7?�O�э�Q��^O�+x�~�}�o�v},V���	��<x��y<��'�Ӻ��1���v~E��W��`��7���w�����]���y�~|O�G�I^����_�� _�o�	}��z��~��T���[[{��S�6q�����׏��T��x���~������xG��ґϳB��~׆������x�K�����};'u�c��޺V׉�+��<z���:�O�����D�U����Y�~���~��5:Tm=|�����qO�_o�C���c���7�xl���ڹ?��+���O��+�����_�G��#Ă�7���F�2��~&�G�O�^�����~�z�i1>����^�ꍾ�q�����g���>���|��p��՜7����R�!�;!��Z{���?{>/E��|�P����qɝ�M�����������������?�l��X\/�/�ó��~���?������m#�m��?xH|��G��z��2r������k�����O1��?q��_ϗݿ����Ǚ?�$�������s4������E׉O�{f���^��х�Ї���~��%߹�V{$��O�﻿����a�+���c���x}E���O׏wi���5�ϣk�����~S򭵉�۟��1���Q?�_����m_�x�?��z�"������:������
|����W���[�ߠ��%���~l��$Vܿި����ŵ�����t�_s��7�����wn��ג�G����#�����5�N|;_��|��g��>O���B���:W��Y|��?"��p�|�|�����ܣj|�R�D��v���`�zk5o�����^�WЧ����o������s�v�}�����U�~�����^}��dr����|~�[���t~>T��,�~Z׉G�K��`���t?�/������$|����^�"�����`���6>=4Ƈ}������r{���Ӯߘ�ߧB����W��]������:|��/���I�x�n�W��_����������K�c{kx��|�x=��y�؞����9����?�J^��<�3B���O������w�d�Z<��gu?���C��������Ւ_��O�/����>��)1�'�8�Fw�?����?o�>��=��������"��n�x��?��������~����_����o�'ޟK>���.Lh}��>�D������������7���g���xwL2���R�ͯ�?�[O�����<���j�#����B^a���f����^�$hL_�:��]�w���������~��������P������~Y����������?�9�T}��b�����_���������h>OdS�?�P�zƓ��5�_O>9&���|�+�8��c���<��|����������nA2�+��٨v? �g|yz��7��?拽��n���[N�����,������1��wƇ/���]�c���X�9]����j�����~�ֿ���F��z��j��w��g]�������v�z�3Ī�3{����p��5>^�}N̗Xt����o����8��_\_�
}�G���p��z���3C?9�����;�^'�y�z�4~j�	�#���]�g���}۾�8��p=ǳ��}|z>ϫ��c�9��z���? 6���{�g�Q�S���=#���!_��?��g��w��U��eο���4���X�τ��~?�����5>ҿp�
��I�w�o��;^O�_|�|����G=u�d�����z����`���\�ګ��1����%���>(��;�A-`�ǳ��ǵ?��g���G�gm�����������u����o8���_~�����+��a������k4��[sؾ�\�o�}���'�������o���'�b����m�σ�\�w�����E|�תݿHm���N<�?I��~ǉ���#�7���5�Pm����C���~ֶ�s>"?�KިO�{��5�w�=j�}��dn����_���y�+�����Զ�;r��b|�'�w8~��'�;�p�|�~�S���X�c�6�� �x*�a�����+�o ��_�e矣���_Пח��z~?�%���FW��۝��Q��z�t?���2w��Qo�/���"�7�S�c>����U7U�=_tf�7�-����o�7�L2xr\�J��1���-�s�d��_�/�����~&��������K��3c�a�Ƕ���W����g�ݮG���-�s��=|���p��w��������c�C_������>`����n!���cv�=���p?�g�{y!���T����<����1�r�ﮖ�p�#������3����	����q�Sa?t�����Ϝ�z��g^U��J�ZZ������x����=,��5��'��j���_�����`��U���H��|�p��l���[�/WIf���^�P������I]g����X5��8������>�I]?Q�y��j���j�k����;b_�[�$��'$�?O��/�k��y�o|e�ޏ�ܽ���ӟ��&���o]���fl�:���3����-܏��^��^��9"�^���e��b�)q�����<)�a�'�~_�a,�'Ğ����F�0�~Q�?}���Ѱ���c��χ{8^�=�7��m=����_���d�z����ڬY���{��1^��K���������v=~�Z~L?������s�_�_yJ�_���񁹸ރ_��|8�C�������5|�x��>����r=��e��?������/�:sq���s�~I;>�z�|4�������?��Η��&��������l�{�dz;�%���~c�����}����?|��{�Z�������7��#�~�7���;�3�W���w�i������w���Ś��5�}��������m_�;}�p��j׫��Ƙ?���m�������ĺ�b���;$�D��^|��g�Z|�����5���}9����m�����������+��|����8>������|�|z�d|��ө�t��s$�Km���������g���{��o�����/�E?������$� ��r���j��;��{�}���u���-����'�x��m�@l��`O�y�����x����^m?��q��|�aɇc|�[n��r�xt�?8&��q����%X�z�����j�ԣ�s�ۋ\���7�z�������r?�|c�����;B�����Z������z�'�W�M��Ca��[�ܖY5�~o�cO��.1߸ޟ�����o^�������7��~�������3��?��'�Y�}>	�1�+��7�]��?�pK�	��~:������_�zZ?��U�σ?8^��g�o��;���w����_�|U������-������w�?��=�_��])�w<����d���O�׮�����j��95�Wh!ܢy�*�5_��_+�a_����SC_�/n��^�3��[�y�`�ף.��!/��������B��O�����z�~�#�'l����o�x��?ğ��~�u��M�Ok�ۿ����_���*��������֧�ۺ~���\\7~^Sm?�;B�ă�_y��u�G��>��<B�7����g{=���������������؋�Ϻ>�wKm�l���˩jϏOΗ������s�s���������
r��K��1��x��'$�^`~D/��a����\?�������<*ם���'���o���~(��7e����x>�b<#x��O��'��������b|p	�7���?_�el�ψ���}�����M��ks���m����|�_�_�g/�:>?C��B�j��̏�f������ɰ��K.�-<q=Fnp���������O�>���χ���q��*��O���cK����+t>�p��\��{;>)�O��_G�h~?q����K&�>��|O������tl�~�~���k/���=�=�j>C�G�C����ßO�x�W���o_{~��)�E��ϳ'\_��ҧ%�U�����	���j����-�=�?����m��C��;�`����qJ2��|�\���k^Oel?(��y�d֒Ħ�	�v�a��޷����������/�l=��ۘ��P�|=&���0�F�K����}ծ?;�����$�U[��ӟ w8�=2��؟ɍ�b�xǳ���j���\��������\ϼ �cO���q�d��	�p{�O@��o�ﺾ�^�s��=�?������~��uGc|�g���x�>}�~�|I}a%_	�r��+���G<� ��z!����ܼ~4��N�>����ߒ��E2���ԋޏ��x>����^3bl�G�Gt~ Ϯ��;b�%�fC2�����ݏ�}���q|�)�,�~v��U#2�����/�����/o��9�����/�z{<�x�|���Ԗ�?�o\)�Z�ﻸ�����F�Į����F���U>{T2Xs���f&�<�/R�x�~������OW[�Pϛ���� Ɍ���U����z�\}�䗆��u:o��W��*���yR2��|L|8��l�#�W��ww��-�?f���m����%�b����?3���ݏ��VNپ�،�ϋ��{�C�s�~I>�U2�)~��W�F2�����q��z��]�j�s����w0���K�R��S��O�ߧ��}A�o�+6_�ގwt���.Z���_��s��W���e�_����j����>@|y��xu� ,t>�x���w�L~�'���>����������
��~s��/�Gp+��=�	׋�9�)���K�^I��~��|ѭ�|��X�|����pL2�����-������B���{9~���\d� ��%����Vm� >�~���7|2����Zm��W�̿^�f���OХ����O������|�����Ч����^/[�~��Q[�> �|^����?����r�Em��%��u���2?�[�Oo���k��{Ώ_�'ߺ���?Ƿ�������'���p�S����\��
����Ķ�m}<�9��~���>��dzQ^��^��������_�e�7�s>|p��a/���U�T���ׅ��Ӓ/����w��|��rm<�|���������t^�4�|���?�g|{�!��~ O�~�X̯�=�߱��H�����d���%���.��� �4����"��O}G<�������a����Ua�S���W-?;\m�=?�Z�!W;�?W-��[�W��oE�/�-�9c7#�8�?�7��a���O�=��`������Zjk�7�Y���e���_�L�Sj]�/�����ϓ��?����6�5�����8��_m?�q<S�(�r<3v�+�t���_����w�U2�������T�>b�|�X�~y���l��=�/���Y�[�������7YK0����@o��C �����k�
t^��k�����O�Km�9���������=�7�{S��w?�j��g�_7~~m؛ZO�CzA���_��x
W�z.�<+��B2�xD���j�~y߯1��Wo������`��$�O�c�=�_�*���B��B���W~���b�J|}dD~\<���Jɬ��< ���*��I�����w��q�d�����C_��珿~�3�����-c��%�/���m��G�������З���7���7�>4��Ϻ��z}��ƶ���D����h��b����^/~�O2�t�%�;����gћp�}{��r��?��ﺿ�?%�v�wrR��:^��W�o�S2��?$S/���|���ţ��e`�����v?�=)�X��U���A-�~�[���p����>��`�� ��NWۿ����j�-�T�w�i�������g�E����������E�;����������l|�9~��^�����q�y>�Do����j�,�~��>�����ĺ�`��c�}*������?�5��-���'��|���K��{�:���G���Yɗ>��m�/�gWH���0�������u�>�x�?��(�k'%�P���=U�~)��H&W���?�$ӛ��>li���j߯v���D��^o���?xh��7ͯ�5����x��k�?��_��q�Q[~^2�%�7 ϯ���8�ӏ5���OX��z���<�:��nro؇���z�}\'�������� ��$�����Uۿa��/�Z���w���7�����/S�������������8���������O�h}��x}��ob��'����O���&���K�O�K?+��j����C��*��V�~��_+��w\2|�x������Z�������o��]]~O�KP?u��ߟ?]-�$VO��\��B�}9�����o��{ݟ#~�o���{z����'��[��c<�_�&���t)|��6��u���5`��%��3��_������$���R��w���_Om��7TS����,����3^�߼R����\c߾�l5�'����1�1�����Z���3�~�;Z���t>��=�o�D���{�>���	����|�i����y������L����8���?`���+�����?�������z���ī񊵓�������׵������
�o������͒�O�o���q�T5��>���u�?P;�����K�55�w�r��Z�'|~�j�o������?�^/�\!��dm5�8_��^�E�^O�����rZr��>����#z>|����s��+��uN�>����������[���C��d|�����ߌ�y<`���p�z�����ϼ���ぇ^�o���?���O~���O��֜����?����8_v�o�3j����5�{_]���۪�ׯj�M��߾��oO޺�����o��J5���t�7��j�������:b���O�?���ß���6����\�ޖ�^�z����\��1�o����h�kR�k�?��T��������'%���7���o�%NH�^!���Ӓ�$��k^��t�9>~$�G>ؐ�w���|$���G�����I�S`�Hf=��^���j���w�y�|��\�����3�S׆���!���i��$����2>ѻ�L����׽_�\�|���F2���ܿ��w��9�V���'~�V�����Z�u�^�K�������j�G'��?O��D���/`����f~�[�p'��?�:ߟ���#2X���~>>���;���q���:&�M��t?�{1�C�~�c�!>�wϮ�wLn���u���߉�[��_�̾���&�N��l��{|h�:�z���1�2�~�����j��i}u����?��o�6��]�#��s��W�?_s�f�:���������x�;Z�d�y&��~��*�'Y�z6��|�jΓL�_t��,���2_��_�{�^/��\��j��$�]�����+������5�x���wC�F�s�^�c�^���v>=���·¾�#��?�r��y����Fz���#���ZI������W-?"w�"��}��*��o��/������~Q��� ?0~�I�Z���}�G����`��H���~�m���W�g ��X��t������ע~g_Ϛ����w����W�~p����~4������O��?�����l�qZ׉���~���3���<x����9��g%O�C=_�z����z��g���:|����������~��6�k�����/�a�3}~�?����H�����gm���zA�+=�����~sr��sr���o��^2\��}�D&?z����|�E��N�m�c���Z{���)��~i�n>M-w���o���z��C�:��&����O�=��/�?ʇ�Ԃޟ�T?��GW���~
W��d��B-zZ�g=I���������~����}?���5�jsσ�������W���-�%����c.�_�P��&Y�?����#լ��Px̔���}�֘���n��B~���N���~�}~����r_��?9I.����j�����S���/$6�Ϙ�V���d��~������}{P�����b��/���/��W��9o��2_+���)|���d�3���r���x�w���j�u���f?%��y������$����ܲ>�}�{ \�c|���j�sP�~'̿��~'s��ޟJ�����B��&w���׋��Xt�����x�/��^�����^ϥ?tR2��w���OU�����p�6׸�?�g�������W?^��=^�~ ^���X�O��������Χ���p�rǗ��
��������V�Ϥ�0b����bB��L��u���31ޏ������3�}�7����������d�@�s&Y�?�Ͽ����O�?���[}��p����������l�J.��������U���x��k����j��WV�����\����-���A,O��x��KZ���o<ŗ�����?����ɫ��W���uܧ�����x=xW�����X>+��Ś��n�W�ow�>�x��A�w�?'B�Ģ�3ה�&��'�����wk�7����(����]���^�s����^���[�۽��cٖo
}ro����0��oT��b,U=���'�价��Տ��[�y��R}��?�#�&x�X����>�����ׯ�k?|���שM��}�@��Z���	�?�^�����?O���x��<��뽷����z�/[{��y�>�ܯ����S�k�$k�ڿ;I-1���>_����z��|>��|�\��?�Ϩn_g���ۺ?~s5�ѧ4��9��드m��Bj��t���=&鍺��j�Mq��2�i=��O�7q�W��L�_�=��<k�Z��������k��F�-�ͷ���L����7W{ޖ������o��M������+ޏ��j���5�ԍ�ُ�}��X���m�9���~��|��������l�o}����4�A�Z�$wL�_����F�?/���|F}`�N.�?�X����v�|��d|����#}?��d�Z��c�������_���/�y>O>/;_n��c�_����yG�]/'�9��/:o6I���W�#<���x�������_I��ߟ�����ֳ��k?p�/:��3v�'��N�|����V�O�Q����q�<��~-�v��|5�j��F��>���r?���������٭~z�9~�v����[x��p~��R��~��۹��>�_����u�bB�?}�o��wu_�\2�ϓ�T?�M�^��߮_�'�Ǯ��=l�������/M�~�x>�����[�ǻ����tX��W갣�m۟���E]�U���N����?�'���Qg��}��W��S�ϧ�y�_�_�w���z��;�3�����������a^�;�;������A���*������e���������$\2λMh=�ǟ�$���K+���߶g����G�|k�_��������^���I�W�U���j<=�Y���~����ϻ>c>�sr�׻�z����������D�O��}=��a�I���?g< ��o������7~v�ܼ���I_z~p]�-t����z�t��s;���y��j��}`����5�k���n���"���o�-ƣ�r����I�U������U{>�P�<�z��~;�r=���?�|��ʮ���9�-w��P=VNz??�u=���G����,p?�g��w�����;|jַ����x����z���o��e�������|s5�-������z'kY׍��SΗ�C�C���|e�?)������G�7���+��Ij����y���i]�,>2��~'x�|�^��5֣���P�?ks�%�֡��$���k'�ǖ�O��{�������u���_��aդ��>���S�o����cw�����`��U�}\�w������囘F�l3����|o�|����t�v��rE��g֪��+b���n�v�X������~H2���������z��+v��P���O����>?[M���W�?���g���S�#gV��p-�ך\	�ӿ6���n��%��x��c|�'������[���kZ���w���{Z2sQ��O���_�9&������q�����j�otY_���?����Jx����B��xw���$�o�3_M?��+e~�?���?�G�&��u�l�O����߽~G���q���A�����/�����-���o�'u|��g�[տ���~�߷��������������|��'��륮��p��_�F�p��{��w���~"|B�K��������M�M��k�=�=W��i[f��񎱫?>�~S��b�FFi�:k{�������֞����>TOM�;�����#g'�o�����������+���#��}���O�M��S�5�����x�M�>����Gr��o@���Y�;�����~����}�����}�_]︱�}<���O�����_4�A�C�/w����~��x�^�ۯ��I?�������ǫ��v>#{u���D�y^��s~_�$X�x��J�_������!|���W�����],�����/��X/4�~C��罞�ڷ���������
{�:�:E.�=/������{V�?qa��پ~e5�b
.b�!�x���"��/����r�7�.�د��|x��-��.ڬ)��Ol�������5��׆�:]M���+Þ���J�7M���������[����<��r?,�~5�n9���';V-!���W��aju��Ɵn�>:_�p����y�ɟh�7Ww�����������ޗ�7�����p<���/�#����o�ݷJf�A�=�w�<$������ٿ��#�D=��j���K��S�^����<�X��X�+z7^�}ޏ�������Ӓ���W`?�%�3�a�7��|�~��=~,j<�P���7?��Z�j�?N����_�_�j�����/
��ŁO�h�c�7Z���~���?NIf���7��A�-w�m�������-_�"7�?A}���-�����ÿ���m�KM������{���O�~��g��硈m�"��/�����j����m5����Z����{D�_�y|���(���!�_�xi���xHן��C��L������=^M}>yS��)�����~��ͺ�ޛ"���'�����,��K������-x������Z_�kx}��~����￢�g�o5�El���m��u�����׍��4������{e��$z'%���Xf�������Ք�=ų�g�'n�>�g�=�����	<��7V��Wy���)�D����|�\�~?{�ܿ����O�v�~&���_�ꈿ81�V�~,|E�xW��U���΄���cg��5��gC�ǫ߳w�������l��_k�>�|l< O�e
l�~�)��1��o��>��~$�[��~��u�KO�,��T���+�.��ߦ����E��~�>?�/��w|������	�a������|���r�׷��ח쏯�zm#����_�į����ΗRϹ��z��/��������T����Z��9��o�����$���(Sp�+t�-��������}*�wh�ǎ���$�����n��������]����~$���j�L~k���8�����<�+���Nh!�o���ڣ�o�~�)t�����~���'X����_�����'��o��u����N��z	?S^���6>�N(O�ޤ�ɓ�����W���L���)�M^?a?��S\S�=���O����;�\->���/?�f=y��^x����)�r����G~*�o�|�����o`���׷�=Eo�����|��~5k������S�
�k��}Ŀ�|���x5�����u���}�:�l���X�/kc�ߟi��ވI��:~8�����	Oh��'&N����������������nh~�ш�׶�`-dR����V���0a���j�)�Y������u�a����޿��h�A�l���Ŀ��O��ַ��5�<{/���o��z}�O����)r�)ɿ���m.e�f���������6O��M�N���U�+�ϏW�����I��F5��z�t<���ռ�����̗E�b���b��O��rӯ��h?�T�/�t��9�+�|M�gf����]�\5�oz��y�N�������ը�9Em���)���g����c�/Lќ������vOx?Rg����}��������_�Ao�]�l��ׅ��Z�y�/T� ?�H�>|�>����M��>o����S��>����������Y�?����?��'�o��l=k�U���b��G��_�u�^��o��|��9i<��������{=�|��Bχ���?����ϳ���b�qJ����_�~���C}��|���j��L�k�g���>����G���O�z�w���k;�)b��U;>=���{O(?q�pR�5�\>'��T�IƷ�?�����P����<��Y���v=��o���}>��js�x�~2���?�v����g#>�����������n���	��~������o���6�| �x���yA�������v�:���(�B��|d�:E���E�W�S'�]�c���N�_��h=��i�O�Bӟ���	�)֣�0E���	������]_�Ƕ���)}�t��~����n�M����l��&����M��	���N����i��)�C�q�#X�t��E>������_P�����"�}~�o7}���9�~�����S�gQ?f�^������6�.��]>����f�s�]�;�����u(��ߴ�W������3��K�����m�������v�}��7����z�~L�_�_]S�g������$���������x>��|
�~�ib���~+��\]�A����)���b���G2�F�S���!���/|^��/�?��H;�'L>*����k����ir��o�/���;-?����.@kӯ�d���h��'��O�{�+�~�xw����f��x��O[��W�	��i��¯>]/�+��f�����K���'�WZ�����T�������w����q��������������������fe�T�Kt3}T׿-����ir�����'������?����\����������]�T�N���Sޝ2u�>km�e[�T5�b?���Ğ��<SGg��/[�����j�3�o��؏���;��o~?�y/�����bmK�7=�����Ex>q�f̞����/to���B�g�z�x���_���m����f�a���Z���Uݟ��Ӯ�2�>NJ�wR������w:o?��Zקğ��v�=��]S����tw��{A]�{/��N�X�2_���z����z|U��^�i�'`}U�y�%��N�~�Ϝb?�ͺ_�+���S�E����ksO�?�~��Z5���[�ο��u����7��W�����?��i�ߟ���o�����>�ԗ�/�6����3��������gS��ݯ��6��ٛ0�zb�k�G��ܠ�Բ�oDo���ռ�e����M���������o_'W��;���]���j���V�z����[��>��C�S��O ���@�?t��~��iW�x?\����uZ����kJ�~?�m�O?�����]����n��;�����������v�p>� ����>��ǃ�v�?)~���6�쇟�����=�ڜ���:�3Eo���R��;������=��i��4���8E���[6��)�M��W~�b}�����r��z�����;c3�O�~5���g�S���h���*�߰��r�/������WT����	퇝&�k��ԯ�x5v��S���3���v���ӟ��g�Ψ��Q;z��T�j����g7s����{�MZ_�i񱯯���?>⣋��������I�?���#��w�|j[���������ֳYOj�m��J}~s?���Z�c}���)�S����8_w󝔿S�N*�����l���Y�^��w���ct3��"����\D�e�����z�﫪��釷������i���ߚv��լwM������}��[�g����{~����O����5��m���h���6���i�b{����ԓ��O8�GլÒ��w������]��&�<��E��o���N�m�Dm�M�m�z���'��ǆ���S?w�޹��q��V���������N=a����|\r����M|�����I�+v6���[�<Coϟg}F�7M��zE�uM?�	��8�\���/MQ?�ߥ��J�����������I폣�~��g�y���VS����4���p���״2��پ����3Ą�}�=��5M��θ��b�:_H�G�s�z�=��T߳��3׻ϺC���_}~4�n�����OS���w�O�:�붰���kQ�������P��:�N}9�z������g����j��f����:<�y������#�ϵ���ɓڏ>���Ԛ^ߟ�_k�����;6����J�r��W�{��Km-��^�t���6^�o�?�s��,��f�����U�g�-���v�췡g~f��_(��/�_����O��N�ߒ����?��ֺM2���+�w����k����[��ޝ��LS5��ir���;}����k�c��D]'vԧ>�C�G�	�W����9��_�\������?E�<������3���3S?�~_V�}�w�z\�e���>�R|x��m�9M�J�z~f}�B5�`�zG��i����o��ѷ�?�?{�w�Qm�3Co���GV߃;s������3�[��������/�|����~F��yF照n�Ϳ����?�����+�w2m��[�7M?�ְ�ֿ�^T��ss]|n�|�|;��j�f>������馟>Q���ݎ�L�?�a��[��&{O�n�1��}R�����#�Vs����i��լ�Nw���CM�'�뿴�?M����~�����X��po��9��ѭ���=�?d��5&u>��`B�U{�?LS_���l�g�׍��S���آ��i��ڟC}9������_��ѻp��m�n��1�ﭦ$_L)�N�^���_~��}�_����������l��4�����8M}">5sq�����ק�����M��z��Λ9������z��ê]� >�?���i���7������~'�=Ӎ�Ob��zS盓�C�gU?`�`m��Nx��ͻm��[�7��ה�_x�>����n���?��v=b#�{W�o��cn��Y�s���V�΀g{�yr����e���>����x�ؙt?��k�۟�hR�����/ �7�p7�)����&�_�g��~i��ӝM�?�k������?*���K��i�=����W|���:9�#�{�>�AN��LK~����k����h�s���o�m_�oR|��qӲ?���9z铪�g�Gj?�g�o9)���_�g;n���k�>�O�;"_v|}�����N*�Lw�wR��w�I�/�_�?������r��yk/3�l������L�k�/a�Ȥ���1?��j�K̼����ɯ��M��u����;��쳃^���3o��ӯU��{R�Og�Rߠ?4����z`��j��;���]��~-���t��y����o9C>����3�?�[|i�z5��f��?�|P�;���g3��x�q϶3s��z�z�G�L���cf�ߩ�������3�O�wW/x=a�����ϼ�ŷ�կ�����M�k�	Xl�G׶OW+y�{�u��g{�����׿�;�mT_��o�~�g�}�;�=Ճ;������~��S�kO;��̙�3�]���3�����Y�������L�����P}���l�/f:�t?`'�D�������]}��ܙ�kO��F?�tď�g�~?�Nr��[����~��_F|}�����t\zBx0��Z�_�a�ق�������xt[�?$~�������i=o�a����-^휫f�Lk�Z_��N�����Q�_ts���x��6����_��6�v���/g�G:_��xܧ�u�7����j��\3��|o5|��������k������\�zs�-��/v|W[��^^옯Ϳq�%�h3F�<��O\��t�����Į��;ɏ�̱j��B��?��-w��4_�jR��fX�?��W�G3�M�7���#��ų~���v�i�zrJ|jǛ�y������;'������N����ow�����;6{�g��>�t���S�_��jC�Of��k6�C����-z>��~���7{&g��~M����.�_v�lJ�#�]lM����P��g:��r���?{<Qo��O��ϼ����3�4�Ŀv�����N���p}�wG������~G�;;�'_uVf��.���`���.��a���SZ������]��2��t5��{�ӕ����)����5�3�ҍ�4~���v��������Y�{k�h��m���g:�r��˧3�O��kF�e��Z��A��|����ۥ�.?������)���|�;�͎����-����u]m��k�:\R�q�_����3��}���O�S�W;�����|Rm�cy[�|��7��o��|��S��Cm=y�C��5�@�ю��ή�W}>f�G�Y��y�f�}��߿�&u��P|�$��_��l���떶�4}�&gu|Mʾ;~�œ�M�{��ig��ﾓ�����t\oZ��X5���E=!�5�_4}�M�<s���ߩ_�}��܍e��l��j�ێ��=�����͞Ι�?�3g������*��;Nh~���g���Η�?t����x?�޳��&�_x�����S|~���]�ge��.��g�Y���3������P��.��{O)��;����|~!�Z�����S�G�����n�����y�]�p~8��N<�<|�
�p�sw�Z��0ْ/���8��?P�N�����_�3�a;����|��zf<�r����'U����!t�����>]��ؾN�@�/v^��&s��]<Oj�~��kPg���T|��7{�g����i壝>L�����j�S���7�|�sbk�l[�vZ�n����;������v}S���ݔ��"�2�~��{?�������/��v��~/o�5�a;O���E�6����u����ϝݿ3G��o�\#<3�o��ag����~�c��p���}�e�X���e�=�3��)=���̿��U_�����i����.랯~���Z�7��T��B��T�\L>U}{��6�ж�K�m�?���ߴ�-X7�|pA�S��v�?��ӵ�.fm\�>�Կ�l{~߹D�����#�aZx�R�ߏs�Tۿ���+:��i[k����%?��ׅ����om���]���ċ�X��j.�l��'7�L�����t��K�#�螧~����_���?��x>^��������Kď.��Ϟ��kwm���=�3�{r;�]����w��ȶ|)���Υ�����V��������;�7�������_BV������:���G=����'mb��?���_���v߹Aׯ���y�7lrv�o����V����/�^\���Ym|^��23ڿ~A�w����y?�,����������R��.�byF��,��[����ة�ǋ:l�Q~��{�N����\�<���w*�.���˙����̙糾�z��uׅ��t�:�|r�o��Q��Γ�޾|�D���w���Ns�y�kK�ا��N�j�%�vx1�z��%}���s7c��K��S?s�.�M��ݩ�����v)��_y~�n�����tm��c{<��w��ީ����_�o����:]���|�v�Lʙ�uX����׿Ts��Ν�{��e~�}�w���5�3�{�f?s�Ë)�3|I���n���|O����Â)�?����˙�w��C��+[=�-���-S�bw7�i��.�����;X/<���Ӫ��N�Y����.P?���|�ϵ��l��;�Gwu|dV�W���埻�t�ۻ����{P�m�~���:>}����u��V�������v�}��g�������N�ϻ�U��'u��6?ߵ�������5��~`���-ߍ���s�O]�ܝ���K�B�t��Cx��{�.��u���>��{(����~�����W�v�޺�����;|�R=u����X߿���=�3���N��'f;,�X����\�{ܶ������];���)=���{6�ej���vw�ʅ����Q������ܭ󕝊��]�u���j-�?����.�g�����t\�z�=>���r���\gԟ��_n��n���m��~�{����p��n�Ӛ�=���S�;���;+��s���=;��)��g����+�,<���^y�n����_��'�x�n~�Oܫ�������x���w��ץ�?�뫻�+�ܧ����_w���C�W�;f4�/���� _D�L�]�~fs˙�w�r����R�ϼO�_����C��=��ә����t��/d��A�_�u\���~�l�̙�wϿ�Ώ����g�y��oO�k��?���W����K~�^'�ÇKe��N��y(����a���}��v��]]|+����۝��/��3����٧���j��ʗt�K���x�D�g�,<yh����K;,������B�w�^����n<ޯ��K���Gt��%�c�|{���=;[=@��C�_���;{�����b�嗨�_�r�����Ξ�>_���OK]}2��2�����?�om�O�[K/�zȳ���>�W����D�{��U=D���=#O�u��!|��˗����?�j�KU���k�C۪�'j���3�{镯 �fk�ާ�~���3�u��?�ʋ�[yi���C^Yؒ/غ����K�/�����/�+���/��c\�_,�_��/..�/Vⱋ�)�c���1������r�b%��7]>�X^�_,�\�W�)+���x���B�"n��Z_Yʛ.��_�
WR�+�����V��'VϘ��m�=p0����p~����r~fa>?��9s`��7�9����R~��R�������3�����y�������|�tia���gΘ��oV�h~y�ky0�|��r~ke%m�2x��Bjl�@�gu`����}�w^��w����I[ؿ??�?�ea���\���BF��Y���́�|ց�����,�>�������Ϭ��oR�K���gv�ɧ/浼?����O_^�Ϭ�������Q��&ǳ�񵰚:<0? s`5��z`~e~�ρ�+�����B�������B����J�����y��Y���u01����7���S������..�,��7=/���(z`)�����K���L��Z^�g-/块3޻��V^���r`e0�Ռ����f��~3��J������7�$��{;�Z�&�9�|p���o�o�ZX��,$�<���f9s`����M����Ą�3�\L�:����ZL.qpi�������./�Y�ge!��2��Jfƃ+��W�����|q~~9���8��jq>�oq���g�3�I�\ܟ�Y\H�,.�>���or^�:��骘�o��.H����>�\tq11��՜�ҁ��R�{������3�l�K+9����n8i���,��D��J�� .2�� EW�X�ܴ������R�&-�4��fiV%�o�[��o,�ψ[ZHOX���Bf��i��c�#�g&F-�pi����c^N��Rn>k9q�s���J���jb������Mb��j��� {v�T�y5G�ф��o�o2v��Gu�9��ɧ/�Ol�
������]!��I�/����)�o�>s`]�����g.���m���b���R�}y)3��Rf���-/%,/��4���D�.-糖���~��Y^�o�$�.��5���W�"[T�]��,�{y��˫��˫{2~W����`�&�pe>Q}e������ʠ��~���98��j�&��ʁD��7��Y[�*��7��$]9�����������U��b�@V3��,��4��RzB��+�Y_�,���8����qeP�X�����+oYId�RJ�y%cye��+�Y���g���fq���Mz������7�7ɚVȿ:`�Yծ�Z�釫��W$���:nu��])��Io�~�#<8�����&C�~��8�݃�A�t%u�k1yKGs<�L�����+��[KY�.Ƴ<����3+M�+����f�qu��,.��M�g���_�ɨguH��j�t�Wg����TXg~�p`�����V�:�gu�M��jq0�+�'X|����S�spi��3~�W���/��,D������|g~��0ǳ%��_-n�������>q��;���
�W�Z�?���`���ۯ'��<P��j��m~JkWgup����v��At?9��g�g���`y0���g~u�(�������mO������~ja0����/�]�:���&��5��+��_���ա�V��Q�|����~��_�_�i/M�0?p���������_���0����Z`ү�hgK�3�:ۃ:���.8y����,>up�Lq�~q~���b.,�|q��@�KCk��,�Ww�����*\^�j8��A<.���0Ǖ�
W�2Hs��Z�~uh��AVXX���� ��}��}��}��ׁ���,�}`�����Z|��@�ݯC=�0�~80���A���e0��+�_-G�4�0��}`iq�Ł,�4�<?����M,`����B+zw�l��̯V<����B�+�V��_Ђ�g�g5@���������_��������A=8���g[g���>8���9x`�r�����v����f����@>�4��K��/��<�_���X^�~yy0�偛\*��. �jp��A=�2���g�Q����@9+Zppu������0������� �u$m��A�,�hbq� �_�P�/���^�x`�E,�5��N�xpx���{��ų;W��jqV�K�ܱ�t��~i�~����4 ���AF^\by�ՕgZ\��ŕA�-�,�����z�����CݯH��� MWѱ4? HK�Z�_J_]2���4��j��������^]Z����yX:8��aմ4,�;tL}u�(gq |K��?[�k��c�~��@d]�7Y� H ��������9����o��a˲DQP��fn�'��$�\������:��6%��L;م	Ed'�Ц�*�r�P�n�;��j��M=��K[�j�y M���� 84�j���_H{k��3����	��LlO-gB�=��� ��bS7�̳1�_'u��rh�:��s }mV�6�C�\/����N�C}��#:�O-[�@D��4F�ѡG��.�����>-�������Tb}ԐcA���6vMR��u86;�`>Ɓx#�@�aO�iA��t�>�������[$T2����75���ʆ�fC#�a�%��y��3�E�}Z���@�"�	-|�=>Z(�I�DN��d�(�s�]�!K-����#4���?��)��̍Q(�F���Vnh
IK`l)����`	������:�=���*�/!�+�Ԅ�J�?t�,���CB.��\t���v��g��ȷB.��]r}B��!!0B��v���~p)��Y�E���(�|؟���;�p�#�@�eNµm���ҕ�� ���W�k��M�%So�Ww!ߕ��|��[��nX(��ChCB>��0r��)��a�؅�-��WN+�	��~_���u���y�(�Ж+�B~>Եy�Gۮ�v�k���:��kV����(LI
�'@�^���W�^K���k!�W���ST��c�㘧��w�����a��P��c�(�'r|u��`J��`|��72�|��yf(�^,s�!_�;��
��8/�=1`����`�{I��U�3VсC!�j�����݋G]�����M��I�e�7_hc��kਡ�t3��+nBlj���g)+�|���Q_{RA�
���'�FtL�ɏ6a�¸�\��@M�LsB��	�nRg��w�Ј�^<B�j'��B�s��΍0����',B~�*�'���������:a�n2��L�Q�-!hB��DG/�+�W����/�(����0L^!cA�\�f���)��S�]p]��[!����|!����Z^��Ы\�L��>��7���"-ī����V=����a`������,l�����Z��vks���V~��x/���ҴF��w��B#8E�x��暶���0{@loδ=��#��}/�½ �b���e�vo����BOl����ۛC�f�j-��!7���r9�	y�a�*�A�������p?i�½Ѱ����N�;���z��s:���~p4�τ49�O��˝�$�?�p6d�$-��=����������`;�=�������v������PO�B<�RF�!� E�

�������9�a�(��x�u6���1��U���p`���O���N�����w���t�C���	!�����s�]ľl~"���#��7"�!���K���^!�$�9���%�\��r������}�N�{"<�'C��<$yR��r�!�ar���
I#or�'\=
����EI��!'��{&$@�9N�I&fG����)��,�㾜�y��B!��A����^�w�x/73��a0��?Q!���\G�\����_h��,4m�S�/�$!���A�x�p!ttE;��(S-�/��5��G�x9�[��j��Ш�" ̎
�r=/�|[3�\��� �Z�(y _N�f(�Z�U��
an7�� D��\q+��n�1G��av48Ciwh���/�. �J��Y��h��q������7���?xǎ8���� ��������4=�|��_�K@�����TN���Bh�􍔐+�Ú>�W���H��f��v�����A�����
���͍�����[�1��\�W����Ȁ1���Р�p��s8"5���r���k�B�RM���gB�c���5�B�
�}���:gc��b�
A��~!,�D�q0!\Pȷ����BPW5�	K���cL��V�B��g�Ĝ��)�]8�ǽ �'bO�0�'�*��H�;��+�°!�ZP�&<���I�
�6<�����(�3}�.�|&���@�-�Aq[$���^03T"\"��B��.;c!W�ִŁ�?!�wkBt,xAޯ�O��[1��i�b�(��r!?�(M�p:/��mQY��.��"����DL����6���ς�r!����c����-�**�+�i����Ҽ�}#���׆�Zsh��H�7
��ވ��6$�ch���Zɡo�c
A���s����vC�d#`E{�}�W`P�؁���P�6�R`0|7R�Ag:��̜a�=֎��B�=C��WZ��8p`r�]!6��Tc��~}�3>��A�v'��3aKBS��k3G�}�"����w�=�ޑ�AB����q�4ĂaGqj���� LV��$&���Cp9��K`P<FGOĀ��Ch��1T1�{���v�amNЈ	�~�`ň��/h|����*xAi�q�����@�����N'��:�xB����M#'�uK��
A�'�i�!:�p�e	A�$�i9��r@�$���G'O2���\Xk ��!'�g����	�����������Q$rc���7��#���[U�H ��7U�g�i�b�@��
- 7���5�>�O�nJ�ʇ�v|.��Pt�|�rݤ����סɔ��Y��N&�,k>���@S!א�̄΁�b�6�?�Y�L!tNp�B-r�[�G�!_(&��*��o�8�,"�U�,^�_~ۓ�|��D�%	��P��ٰ�r�8�'�k����Y̀�.��M��͆�b2,Oȷͅx{v!��
�s ު�M�o�l�}�(o!_ʵ�f��d��@�w��#r%p6�re^����������yNyV�.y�?�tm���R>;R���50V;��Au�ΎB���n"�מX�;��١l���/cgG���0�%B~G�� T�*��{��iv����w$��9y���䑤V�����Cd�>1�]�7��IC���w�Edd�c��r��!7���5j�4�!:������h1!,^s"�tNʯI}�Vi"�i�f�_"�/����0 &l�Јek"k�F�ɢ��|�Ny��=N���Up�����,B��ǭZ�����a1�Ǐ&���Ll��z&��¹��J��U�=#����QL��	a�-���4�k/��..�kB�^��3yWu���A�pA!h��pB��.�����bh�A^��+�������~2�o.L!���a�XT,���X����)}7���Fjw�`6��Hr��M�����$��±�4�=��U{��f!��)u�ސћۇ�B�h��
aS��0)������E�o#�����dt�d��y��A|��胄@�P�xY�=Z�s�)��A�!L�7�y�*��F���o�y�|9��Sk�^h������.�{Q8!����C�ʁ�f�G�rZd����$�U
����"�y��gs�!~��C�T��uft��',3hn��ӓ�z��O\X��73�YI*�Dx�H�ħ��'RR1م�Y	�q�2��I�~�X�+r"*�
/��B��p/�]��w�Dz!�W��|�ԭ���qR&��<�	m��(����Y}��zn~��r2>M�>9
��3i��3O��`�!��?Z�W�VY�?�*�mWU���	"S@.��-��	��S(u_2��kkk퓯�5�Ʒx�88�0r1$�k�_h��&��Qȕ�B�h���%@��!7�B�a:/�F���_���1�Ϫ����Un!|G�r!��]B.DySy,�x,V��ڌԫ4Hh"7
��]�P�F���c��.`�=W�!�HB�!��0�����U)����ځ�h03��=�j�f��p�[.���H��x>Tȇ\G!�����H�:"�
�b,�N���Yn�������C��.�B�Qtu�B����#�B��# cu�D(�.ık!��f��������QLA�=�����W�ص�k���"�����00�O��|ǺvMk �C�:8;|�
�p�]�ӊ�����(��w���Ak G��%Y����Ʌ�9��Q�Ȁ�f��B#8���278;�eB�p�x�Vy����n�p�F����r�Ⱦ�R-
aM��;\%���&g�D:�UN[@�﨓�B�BOL$�^LDZ�ƀP�A�w��N�00�^8��~��˰�Bh�����8!^L1ZME�Q)Q�
a�ͅ���̫6����X��&�wB~.�J�!½Zȇɂ�@���_�`!���vs���� Օ�D���E=z!Ɋִ#�����]��fe=�=��h�aODe!l<gǂ#g��^H�"���n��}l0��������o�^���4� ��D[�>&6�����V��ϰPl��6��F�Bh"����l�WָD��3_5(��e����!�9rvBloX��7��d%ZLsYȟx��\���^�s>!l2x�'�/t(������� �EeF� e����$	&(	�J|񇘵�|�8 P�`���*c�
���@F�-5OD��B�}�sp4�$'���f&M!h�"-�ж��B�/u��Dp����@����3������-c�j�$�!(�.K�#P�]�i �x��ES	*�YPCf�L!~��Qm}y �I��@��4�q�x��\�BPﲡ������B�9I�FҶ��b�Q�O�#��P9�c���J�h
�t+QN������p/�v!�oO='�,�'��[�]��'P8����>�Ǆ#z9�Y����JB�uy���;
��y�)m�M[Z�v�책�TX��ћ�7��7NX�|*�^��e^�EGU
�;�`|?�e�?-ԕ�����Z �wD���� �nnϣ�B�������k��+Lyh⇈����Yu�B��֎���!�_��*耫��y�'�v��&����{v��F/�Ky��A�#{�fb�͔������v_w�u�;%SǱ�fЗ�������vG��2�*��)䟶#jF]�Q��M��h*<#6��m�B�"N!�~c�tԚ�5�������^�����1�'�ֱ�����ԭ��y��wB~��yĶB+��ek3��o<�|#U��ӎ��<�{ ��_��w Q�~P��(���=P�E�p ��p��9o�@�����qHU���HpSux�9>�/2L�\s�f�B�_y�6X�	]!,�E�0�'N�+���ĄG����n����)��H!�IWH�DUJB�\�b9�z�Q�ԁBXt���W����;�G�?Įi�_8~�<����D
5!�=2����֭���ZH�*�q/�Ă�q����/�����N���Cdj��c!prk�M�8rx�UY��C��e�w���B|"�p�B���T��KB�0<2�P�����c}!,��"m��J!���B��6�w��������XK�#���_!������v!���TN7J�T�6&<������o�ms`nD�oe	A��]0����lΎͩ�a�b�x��w�AF(!��B�VZM��Y��>�7�P��)����D�0E�|��ȋ!9qPYhMT�Q�*�3�P�)W�v
a;8�װ��:M��_��%�A(�t�x s@�@&��7P�B=p��c��|����B
a�FǄ	�WJ�@�ƀ􍁕/Puz�L�D s��kBb�8	A��s��z�]�]HİY6nh��C
�@���l��>�BO$oO�k ޽��+����7"�Q1��ډ$dB~�S��ţ�*U�F �W3� �	�����H��H�x/��ڑ(d!��6���R;��X;�GBX2�`2��fm"�xg���H㥭"�	��gn]�8���Ie��U�0y7W��@.��p�Z�?��@���RoB>��>�΃Z�B���U��e���Y%�B.}!~G�9R�
��(��b|	��BO4d��I�h�4r5�4D�^H]s�L�p/�e
�5���j_%4+�:�s�B�����D�4��
�j}x"UU��CX�7/��ډ���v����i��m�,B��W>!�6�#Wb{�"�aKy]W�?p{�.��r�L�wM��%��߫C�?�$'I�q|z�UTMe<�a<���k+�U�f�J��'B�/ī|�t:��Z�1;j�
AtXA2udC=9#*�:�����G�D!�p[���1?�p{8e�ˣ�f�B�9%B�X�N���u!o*E���l!|�����@4��oX�0a���	񇈛+�B��at��耧�a�\U�@#p�}$W��x�6,�B�zk�/�68���~p�N�ډm��Ȑ+��3����*�6"�huX
�ȪV��>���Rȭ+����P���D*�_�a2�S�<Q�,�@�D'R��UT�&�#�DHQ!��t�D����:!�
�;"yU!�6�B�!T�	s�D�������
��o����g� �Y��,zW��q�&�Y�vp*��k|텔gM�6!w7��]ߑ������g��Q�`J)���Vw���YT�O���g!�Y�P 5j%vs~��1����$���~Ñ�0����F�B�
z���\;6*�Abn�����s�B�/N��
��Ms{/�s6���E+W!^K����Q���f!�c`��8:,zwvb�ۨp��E���t�xz� 	l!\�m�Ar�s�JTGs�=j͜CC�TQ^����JrB�L�\��q�IHJMM" ��Bx"U�CQ{�<�"����p�x��R�I�C������|yyW�X��Xx*f������9/����
�.�@�����l��h��������X�B�����*�E;y Z_�_��B�'A�
dЪcw�>�*R�| >�BXE���d��&e���9�;�D��Bh7��@f!�Wrg�<���G�-!LѤ�"9V����{-�Q���'7�I#�4'�����V�D�D�BȜD�	!��D��GN@K���:�������2{U%ԧh⬩b�'��x��\WQ8�㾐wN!��O���s�\.�A������`ňg���[��̢)�_;X���oe!7����O�67T�g_�0L�H����
��r�$䚂^�uW��ArB��
�Ji+.�4�}��s����	��*�^����ը`���o�qB�Z��$:��\M�v�~��K��c�#�ЭBn��M�&rG��`��Bh=TёGDJ��QBLi
��#[ڰ/��H2\��X툥����Ux���"�StX�
���Qء�
A��x��0L�܀�d��	�l��Ql�p/RB#P3H��N!�o�\|�
�]p/�w��9�bi1��:��Q���0��?�*��OK�:`���U��ȔP�_�'j���ԟ8���j��'�*��j[�{A7���N�v"LC�wMUP�B� i�n�r���c��q��iU�G�||0�L��g�B�
i���N$"�T+��s.�CP0M���<�oc�|i,���E��*ke#��YHx�����Q�ĂJ�<BO�-<2�
�s�?Z�vq�.�a�.T�����$c!gW0d���Z��Q<'6Gᆁ=x�#�����H��q�p/��ڱ���C{ܨq<�~[+&n���0	A������F�R!�n\e���F�[eTL�#�c����QȢ
�*lEX���
#��N9!<�����B�B�f��]ӡp�Y��А
��̾X��YS!���M���wX���	A�?�=
�s(�����w��z���J�2����#,:A{a��]�I M�D��
�*�A����O�
����Wl�wa��=�*�~81|)"��b0�Dm�4��-IQ��$H��]���!;���@��S��$PaE�_�֨�oT0�LJ`�#[�hR�MԷ
�B���-}"��9�v�@f�Z�b[$R�	aS&�����}R�H��G�J�(`,�.��΅A�H�+�9��$�0����ԛ�o"¾�b|!m� ����\����V��%�*YM����\N�U�S"��Ʉ���M�~ì�w��Kr!��u،w�E7y���'��BT��t!7�UZX|!���c����\l�;�V������|�o�$V9LPV��	!�B��%#��A�u!�5e�~�<�r�S�?��[s��˜l��	aZ5�O�IJ�!�Z�O!�܅�`,��А�)7'���� �vἣ�Kse5��ݐ�%�W�c4Yղ$fȅ\t4$5-�45|}�&����;2K�"]Ȼ���_ȕi+�	a���������:�G'Oݤ�;��'�PJw������UV�?�-��4�.���3!�Y%E
�^P1�@Xu�:ru8;�������s��@Rf����Gôb�d���{�<<ro����GB���B�!�~p)�R�ھ�b��� !:�)d��������c@�ȡW�������X,�(��0�&lȅ�sL�da�e4!�Q��p&��=�Ʉɢ�w4��ʍ�?�P�H!��1�_�<竍!�EI>�_�<�+��"�D!4n\���A>�O.Edr�Mj�Iۄ����0���T�_HL�L�,ī|�*�և���8
��B�51-U�;y!^妧���@�hl�L[8�I�R
���#r��`�)#�3!,'B���P#YoN��*!�WqZ51�z�V6#�ſ
ᵑC��2�P{�n��D��Ch��B�
�H忌��T+�4�i��q�Zy�Ѕ	�j��|�ɀ;!�~s�U- L��|���ƫRP�^0��ިBZ�{b����̍��B�H��p0r;fn��
񵑑 7�non~*��#8d��j�>���j�أ����FЪ�+��os?�����K�x�..`	5�p'Ͱ�<��.:�f�õ��{B�ۇZ�A�S�������Or{!4�|y�๐_}^�F��/�p�w�n!^�����D�W7��A�!���l�Y��D�!F�AtJ�CP,�'"�6r�B�p�_ƃ(�S��C䖩�G�9����	
x�y\j��Bͳ,�[ �k@��k�0νBPD�\��D�
ac�����U�=a���dp������� b#��,A�b�?e�ƥ�@�Ln���D��*��OL8�g�8B�L���AsgfՊX���8����+r"�7Y0�6�DA�d�d6�Bx"�{�p�(>��c���N�H�9ͼ�v��ߨ=��h{�C��/��>���x��o�o��X�`��k���b�Y�b���łm�5�.��^�-׿����u�����}uO�/���/�����3ؖ���k�k\l�n����ߍɽ�Fm\_��=b�~�<������b�gܜ|/������xFX�/�����vs+\vE�%�x���_l�~�r���6����:~1~�68��u`z��>��W�į/vؖE���n��>�wO�_���u��b�������m�r�ݸ�7���r����88��->��c(?���R|���[���������?���L��o�� /�qگ��q�������k�z3�垅��2(���1~�>�}����2�Oʵ>?�jq����U��>��m��cS��������ܻ�x3��=)z����G�ǘ������ߌύ�w���=?� )�zR����7>�S1<c<|�W��[|F�<��`4������)#��x��S|1��cP֍�y4&���X����㹓:͘�6)_�u�}��g,ʍ�?~�)O�5����q�^�1/���=n��:=�rw�D���ro0��>9n���e>���c���6��/7��l���ٹǙ�z�������c|nʈ�9g���`��6ߐ��~���f��?��^�ϸg�%u���O�o_�&_��i=���QƮ���b\gV�:�>���9�V��n����ߠ�X��e�ߘ�_�������e����u���q�|�w����B���pƯg�V��+���|�w�?o7��6~�,R�v�~{�sܳ�[�u�uhx���uޮ���h|��������~���on�W���Ý[���uw3��F7��q�����{^���$����@'�V�]���^�JZ���N�jR�U1vݺ֗W���m���O�&����pץ�^��R��we����+)���;GH�xM��1a��1_�O�׊Eqq>��	^������i8�����o��W�ǌ˾9��Mp�j|�����P�禗�ssW�&�����09a�u�y��a�k��O�����7��D��k��l�x��y�]_Mj2D��p�Gej�Ho��^�>��5���I���ǺY�Q�c�Q�+;��x��y=}��[�|��*��z�����Ƨ����񵾷���d����y����Mxu�����-a��K�����KX��g��7ʏ��l�L��3)X���Sy"٤��M �WH���(.z���=o��sIN�W�����!��Fܽ�#�Qi����*D���N����>Gr0�26}�ߨ��?o�����1a�{���FJ�FȤ�*m���/�E
���_�^�T��Mg�H����
Um�)~{n�\��j��<?�vi�}�����x�-��6��IгIkR�/�k�]����?6#�|�65>�F���+���5��`��:� ���g���ϗ"q8������`���I�~|�W����ǃb��=�`U��r�u�z�/MU��mW?���9B$�>�׽?>GEipԝ��������𼪕��'Be���|�_=�����+?eȇr�>����������%n���ǩ���K�f }�Ϗ�����C��3�!�c���������"k?�������j#���=_*��g>������V~����|}���½��2��s���+�����q�b�ziP����5�ܿW��!��Ǡ]_��}����!i��rҲ}����Ԩ��o>���!���;������,���{�|��*��X�3��j�z���o��A����!{�|h�����Tk9�g�`��6ۇ9>lm�2��C��aO���>^B`r����"��L�ׇ���>����Kڂ~��χ��ھ6�__�c����kw������_3��r¶�����p��2��������s����ߓ��?��u�l��/��kz��M�?�����_�������L�?`?�î�v�?����M���,뱻/���?����w��{̏���ɸK���;�>��Y�~���I�����#��sk��H��ßu��~��>�oq���o��#wo|��^���ޞCr�Y7����~��{]�?����F��?��'�����c��Ă?��}����׫�o��>���}�8��X�G���3�/�������B�#�ﳗ�����#��{?����G|v����NLz��9��ح��y��������_g���t�ѽ=cc�qc�/��,�qSW���#|l�j���g��O�G|�Ȅq�*��K�Wf�?r�D?�v���q�6��|vw�sGjd:�}��N|����g��s�>�G˜.��k��w_�^̅�`l��u�G�>z�-<�#���9_�!/o�?���/H��}�~e��oς�]�g��z���gm_��vI�0w��Y���?���u��p��J��#��l�Z�qI��M�;�f��Ӎٴ����}���g��z���fߌd���םW
�K���R}c��{F�G���}Ϝ~������<.I���vn��?M�t�M���7O���b��
M�#���W	��yz���'��W��=����ϸ�W�?$Ӹ�@?�3.��yD�Ⱥh>£����|����=?�#�}��X@��pIõ�x����e�	q����_m_e�
�?�M܉ϝH�ݑ��طxY�/9N:��b�A��. 1Z�����{v��	)�Xa�=�����O��M��G����H��{��x�ti���N.���\.�r��ʍ�߾R�x{02󸾚�G]���z�?�kJ^3ُ�\��U/�7����o�����u�<@{�������h�`�Xu����g�(7l �%)4u{����"O�Q�J�
	dm"45����/�)(ZC͈���]��B�hĵ�y���Ԝ@?���u|ǆDN���ä!a�Z���P��V	4
����km{2�r�EO �YUdBQ�B>�^^�y��Bx��̍UWq�uTp�d��XN�H��:�ra����Ó
a���y��-�?����:�#
y�֑���y֓�
߻S�'��x�9��������@�6!��@U�6�'�Ps<qx�N!,cb9�5�]�st�1��B��X�3���A#�'{�B���UD�'�<���}�� i��ʷ�_{>�}Krb6��y�cO��X������3S�<�w��w��J��i"w��0�&ҜB#F��6w�!����CB���p��y0L��*���BXEgz
���^YM�_h!�Pb�-*��c`..�5o�2����B�ik񵷧s���Pj/�E�i��0��sa0-d̒j�ɪ�;�M9�LQ!ܫy��B�!
�7��l��(���$��X���,}B�lT��`��<��<��`|m����B� �Ã<dB��ir��K彠���!wP��|�/B��ar���|���PM?�Y,1tPe����Tr����z�yh�s
A��Դ�T���|���M#�_(�"S��|�Hh|̙W{G�~����"�+��0����.LZ5�[�b�v��|�䪍eτ<9��5��I�Zn�����ҁ-i�H3�?���H�/].9Q,GK@��zm2���i�!���Ɂ\%�Ҁ��Jm _�{eU b뱇����H�B��v�{����QA�%y�����|M+���9,��rI����Ig5.!C���YA��x��{As/����P����P�M�i�w� �7WW:KIu�*�"����#�n����(/�B�B;�B�7��s:r!�k{^������Vo� !_��0ȅ| t�wB��y��w�@�H!̡���6�}`�-�9`�B�jYB#�����$���`奊���h�KxG�ZRP�
�(�%䊈��'�|�����:���O�+�O� �4yS''�~�L�����B}.|ǹ��;0�vי�0�'�Pv�ԩ8W��z\����k�=�$�j^lB��}w-Mj�����\��C���~}�Ck���V����Crb���i]鴛�(�W~��hT}� ��:H�F�.]��QlB���|�ݫ�hD`}��o���ƽ`8�Rs|�nlX� '6��}0�v�e��0k����@B�w���%Y���:(�T���V�B�=r���N��T��B��`n�\�.��>�V!�_�`�"t֌�*6�5P�{":t��P�e�z`;�Y���S� h��"�hW���'�U�x���0�W���%�Up�\�^�����OT_,䝣G�v,	b��h�\N�����ha��J��C8��Ҕ�W
�u0���{��&Lu��B(c/什*1K�z�x`CΤmG�e�x�d�ʑ��x�,*_ۡ�Bt<�pƄ��(4R}*��,?*��Q����9��N!�W�'j\/�ݺ�|�(�R�m�kiB���~}b4r!�v�=Z������;�������7��]ޏ�Z��׬�OwUm�ш���Q[yt��e��&����xō]�wDɹ�Q�]�Ŷ�D�����m|�4B��EM�@���ʟ�C(,!:8 N�*ي�~@9BG����J��{-��2B���i!��c�������*��u !́R�B�w��|���.�ƈ1�q6_���\_{?���u�+qnϥi.?�r7�BhĆ4�ۏ�;�z�P�2m�P��6X[Y���oԘ	Y8��#}/Z~c~��ЮE�d�pv,�4����b�c� �X,�k�E��i�X���`�.�'Dڢ�]��6<+Z?�+��	�n�9>�7jm������§�0dA����82*�n�k�`I��b���Pj6Nb����<BP�X�u��D:��C�HB��U���P�Ճ��A{���p!��31�h��B��S!�G�s�6TΤx�q��`!R!���ZpP�Q
�"'� *�	spP"�;|!��!L��c�\������X>��a������F�DL,`�J�B��܋G~�� }���n�¸����0rbC�	�X�;րg��;�VA� ������w̆ϑ0G
a�Ɂ��3�#"�q�(�Z�G�Ċ�I��ey�{�d�[Ri��-�B�w�	�F��r�s>8����K��Q�v>�
B>|��D8U��Io��G�K�����߫=.�gÖR�
:��{m���l�ţ�+��D��T ~8}{*�ˉVZ�>�f�n��UT�W��`/��?Z�����C����s��x@�ա�
��S�B<L!^�FL�ѳ��bv����t~vδ��C��!W��b^���9;".����x�W���I��k��J>��0�
�'Fw�z�64spLh��g�T�p� ��UB쇎�(�&Z�
H��r�$�ֻ����������Ķf���ʜ��1�����5�Є�v��מ�/�sc���[�9��Os����*��C��>�ɴ(�#�{��� ���5|�1<y�0V6x�p{�r���w��e�^)s��p���^�Q���m~W}6o׆S��������	i�J�s���=�܁A��W���觧�B��~�B��c!����N��>�N�?��?�gb|�d�Q��D*ޑ�/���!�i���������ܜ��� �[�M}�[x!���=�kk����p$��e �ks?8�r���I�C��v���Ɂw<��r�G!<�S4�YgmP�q�?_�{.�f%�v%DZ$v������(�b&�F/�e.�I��d����(�",����[ ��H�UN��a�'�B���ę�L����<$��nO�<ӥ�_*qa#���/M�#�b�!�b����p���\�ɸj�NZ�u�B��r���
��R�-���r�C�v�����)Aȿ�����$C]|��\NH]ŧm��j�J$���ՠv��� Z�X����]��&�rb5��V����\��x"f�b,ҪxAC{!�&�c��ӭ�h��D.��Շ�����rU����p������BG~��-Vȿc9��^���:���p	r�k1O��z���W+m��9��t�j�膍5p�[���E!��c�:�ʝ��2�8�у�F�Jx�}?�Q�,�����Lԋ�2�췎��V�W�kO���������LkB��"ih�#������8+_��֢�p��u���8B��Z�:��
��b,x�WuE���R!�����V���[��vZ01 vs�V�w҅��7�Ԩ#����F �bl͢����7�~�޾�����X6х�BH�h��ڱ�Y^IhR�,:�a0m�ǝ��_�AS_�|/� h|�-��o<���C]���]]x�9Nu.��XX�����I̎������@��Jq��7��
8-7^�i�#�\m+���^���(ɲ���xBG��r£��X
��쑵��	S�b΢aC�6qn� S���pH%�a"��o6!H&�]� ����x��%|�V"o�ԕD8W!4q�B�UxQ�;nf����4��B�����<�*�:�k_e*�헫����"�N�3ý�%䲰�u|��U���||B�FՑ�߾��Yȍ��|w��z�Ud뇆ǺU�o}�����v�G�0�����ﷅ|���ߊ��U>�Ky���}�@�Y=�0V".w�����E����e�iJ�tArekwn�J�{a���v�=rɴ;�B��o�6�2��d�0;:\�w߮�쎸�B��_���i��Q�4�a��[Z!o���8����݈����^A�w�{��r�8�0&fǀ�m!���P�73��﹜�!,�#z�7��<������{`� ��#�.OaGػ���O�#�k���w"wQ!�I��o��+���D$��Lp#�ʼ6�~ү>ۅ^�"��5��f`�2�I#z��2�z���k7c��0r#��r��)�����ڦˎ��o����p���߷����V�؅0Zn�
.7�i���,�Q�����*ԍd4Ȅ��/$�����.K����O�����ѕ���ksӲ@�o#?�fF�B��{bDo����{sw���i��
�* ���a/�{�F}o���ڱ�l.B��q�B����B�iYc����E�C��W���8���N��TD�/�dBX��]!��� ���q�/�e���j3*K+�v�bR�
�^\���v �F���np��H��1�8B�1i	,k7���x@�$6�W ^t�{���?6���00#0 %�� '"�ҩJ�P6|��i�ND�n�B&�¤z�H+��މ�_BXEn�;�$R��<n�>�p�9�p�|������T8� B>r��)�},�B�s�t��:��o��t�b(�b!\�4�B�<B#� �Q �AT�y`��*�ӽ�߫a}<���p��G+�/���?�@>�B��6���@sAOC`!_;N[����Bx"$�F��OD"�B�
��a�
�V[������>r��2u��W�WoW��r��/Bnq;��B�
�@����ӱu�T�w�}G!^��]:���I?<�V=0�:Re��f!ߎ�kB����>�٪����<n�%�*�&�rc��h��"BS���0��0��a|�>�@�)�v�����Bh��B�	DR	��q_Q�@X��-n�ɢk'��ȴw&�`MbU�?�g�a�"!��|�$��d":E��۬�D�Em� �'L�B�V�f=r>HB��'�'���e{�,����_�d!��nO�!k�զ����͏��lU���z�����g��D9���8�<�C�����=1�<�����[����+Uq�@�|�Ю��|���lꫵor��Ɨ�w!�Q;�4��=Rk}�x�Ҷu�4�s����P]9��:�@!��ه1x���|���ace����Z��&��r�����hx�������?l;�j!��̌#�r5zN�[F-���2ǝ��`>���Wu�>���$rlT�#� 9 rB7I��-B����B���c/�&�D'�#���T�B~#���}Q�{B���B!iA�H<Ce�$�-����x0��q`Bl*J�	���G���.>�A�`��B���A���ϡ`�t!Wa��R񄏉�)�F�7*��'Κ��@�k3���O!�Pաr�!y얭h�g4FDC�P0Er4��D��uU%���]��q����8�BU�' !�Q�/���Bh=������U�*��ȉ~\��m`!�v��f��8c��p�B~�J��q?��,;�mF��yZ쇄�il�1&F���S��
��Р,ȡg��R�1:43B#�������{� D綔4����M��d�*� W�9s`�N����Y@0q9���p�rէR4�0�����A�c�'�P
a�O욂�g1��O�|"�A,A�-��v-N��bBxG�H�.��_\E�%��Y\k+����2څr���4Ǣ��8�".�]��G��n��Q�_hs �9���47'���Q�A�膳W0�Mk)A�o��M��QH��1&6Nk� �$��}j���c#qE$�½�axߗ���t�P9��8c��|�B艃�q`{�:
8�K�8@U7B��}`��`��8p���(�X�{5��&.ī0��p{ĨG =u�W �Z����B�
��������M�.�x��*�+�9\~��B��~i�cBqK��	a`f�"�8cB�&��B���9L!4��!�Y	��r�^�8�VѤJ�HY.������%��o��2��U�!�������|0I�vi��r)'��Q�{"��X{r7��t��9�cC��D!��'��W>��5���jCUͤ�����5](��Y��j�gJ����J������\�9rU��UHzT���D$�̄�.����ёK�\���B~�����T?%q�y�|�'��U!�/:����K�/��5	r_��0a��R�@��d��hGu��q������� O�?y!�	�W�F4��C�ܞ�����IcW!^�F H.������%�|#���.8b�4���&��J.'c@�X��0�ʬ�G�6_����_Bi��Bhb����&�0�P���F�串|cP����t��X��y-'���ј�Z���|�X���64�3̉���8��
3��,Y�+'��3U}Gl�JM��|����@!t�BI�\��M��.e�_{�0H�ٹ`�E!trY�B�@.��
�]�_M:	�BB !�V��	᪍MY��%���F����5%S]�m����J�gs��#7B���HWT������w�J���:�ɨ͜��p?t������x/���U�46�v�;�Pq;(��+��A�F!��
�IF���7f����!"���p���͵�6���;��Z�c�J�?�o�;ƃ��vE�G��itb�y�,/����(�}Z��wh=Ǆ��S�Jd�I	�~�8P��Bغ1���@���hMf��D��,+	4�&�
�'�ֻL$�B�'�DJ
!�m�>��𙨞�3�DF�Ld}O&����@Of�Nf��DVar���������Im������u���uW|��Ly��u�'/����I�K>��K]vs{���s�G��O�M���x�������`��n@�%�}���X緼G�?��G���e���T�f�m4��+��qڮ3ˋ�y.�i�5�^�c��[������s7燆=�qӕ���3n��ˮ�����fh�t=����f�x3��w�i�W�'�7����kx1��~#:ތϽ��/�պ_��~�������x��oك���v�ǜ�v�g���{������r\W�K����󸾈/v>X�~cc�2/�1N��|�P�����_�8�Ƣl�^�b�qk/^vV���8���pn��2��r\��7��e��e/߹˒��|('���<��ەc�T�J�N;;eļ�ƗM����#�M��b\��\���rn�yss�MY27��<�;��/'�����=�:�z&�WuD�8�V�\]��>�-�_纵�KɋM��v���������In/߃�	�_?��?X}��s��Ȼp�0�{�v=�^M��P^���������z��n�.�{����h�ו׽���I��&�~]y�ܯ+���C�=���W��[�.��R�|�~�N�>��s�W��f��o��k5=�N��̻G{���|5��Sx��no^�t��/w����z���͍ {7����*[�wn��y�n�7ڜ��r����>|���I���{q��*��z��\�ޛ#�U���!����Yw/}�4~�����%P|����~��1l�3��2n��ה�AqӍ��G�*C{~I�͉��������_.>`�l��/�Wޤ���П�)?���|ɥ���5ln����?����2������|��+}���;)C^�b.lk�6"���2�7��K.]����>��8��%??:��Iy-�7$���{���O��D:�����쓃V�s�훙�5�?�sn�������+F���ɑ��j��y>�|�P���C5jIݦ�M_�����𞽷���4J�򭢴y�ꥇ<*�l�.j�ϧ����t6~g����k�NU��~M���ɏ��5�_��k ����P�}����?S⟿�?�����������ܣ�?��J��ߪ���2��M�O����W�������{���eo���[������޴�?`W�_q���^Oۛ��������H���%�Iǯ~'��l'��}�?r7�?�p�o�d���o��?��^7�G��iǝo1�I��@o�m��>ߏ�?��($��o���&�9����#荍��5^~�נ��*K�nTd���a�?�p���
��'��Y������k��,�a:�^���]��s�����O�i_~�����>|����L��D{nZ�?r���{�������u}�h�7d�o���12{LVL�O��7����x���>�?�z��C��w~��{��#.�_G?r�Yݿŀ��%���rlL��q�3d�h�G�X齱}����]��e�)k/�;�z�Ӽ��W�q|�����R�G�W��|�t�4�W�q���!�����,'�c���;���p��=����#����	9�� ���;�T�?�cc���s����&qI;1��5J���*�G\ӛ�#s�I��m��Џt����GЫ�p�?d=�ut�����^5k�H�ٽn��K�����%�ƿ����k���M�pɶ��$k�>}8]���+ѺN?��Xx���_.��1��k�k�
��,H�W�����⯛��G|�]�%�
�_+Ы�o�.!W��i�"7?�wO�v�s��]��Lُ����
"�_����{�`��c��Z���^-����_p�q{����r�t��1�tI�!����jc��rlo����1���hu;\�y�7���v�>w��k ���������zqnQ���u��:�G��ߧ��u�ϸ���w��u ���{�k"����`G���.t�|E��ʿ�#>���	�8� �U��uK��'����c������	X�le������X��_y�dݫ��4~���#ÿNe�22}����C%��5�^7c�%~�rM�29q)��U���c,6����_�/m��[�ϯH���J1����%v�l�Ye����R+�k}S6�f��Ebo���f��m��}ǚ��{�R��b���#>�r�,H��yM�?�^.�ʯh��[,���w�n}���ܮo�qْ�
*,̉k)	� ��f`$�˟������?�V�
c � �r�������E�X��DMSn���o��a�����J�!=��s��6fZ)�Z<Y��h����P��h�+^5h
��c.��Bs�d�*D���ʅ�H4+�o��/��G�}$�!v��c�<�U$��f5f�iEZC|Xk_�!W���L� g!,ӭ<���꘵�
�<������y�p{T��_�����H��Hթ5�X�I�SU�ylq{���n�!MXک5D�½=)��	Ʒ��	BbW9������pB̴�����Ŵ=�wL����s�����}�����6�'N��<�S��ͅ</E������!�{m���
ᇇ����B�����TF�X�B�/T�mL�#m�#Ʌ0:���'���x<�A%]����X�x���ذ�d���WO�Ә[b�W���~�~�$-�!�Bcy��?����;W�?X~�4&��;"-z�~��a�=P��d�j�hDb�b&!��������.�t��U�_h����� ��<�v�bR}LL����AbNTr��z���q.H��٫f"����+��@	��r��!�F��8�SUa�.\���nKL�^������out��o�\����8m!sn���!��R�mMv����)�K7E#�hC��ژV�s!�����BX���I��,����u�v.�h����k'���Iӄ�4���.§�Hs$��pS��p7H����F�6!6N�с����ۨ$Q�Q��ѫT�7JN���F��Bx���(�^?�&�?��(�)�wDV�B�%�ϡ"�����n�p�v����B�����-��Pi>�s�� ߵ���q:_���A��B�_��a�|&���S� IS;�?D�|!,`gA�;��\qg�h�gsLlL�C�Pޟ���	��*�w;�C�ġ}"h�B%�|�;'X(��O���ݢAtj7�h�|ĭja�TӃf�@M!|�A�^P
���v���rLa�Xޱ2��*d�j��i �ed-.?x�XА\����ks/��-�e.���E��"CZK�,��f�aRgJ����<�!��
A�I%J���0��L���ɦ"�jKIrAt�bS7���
'BVL����*BO���	ش�bn'r�GVT��45��IT��i�������=������g���ؿ���V���|���v=Z��Q��K��	!�k�(��w
�NG�%f���/�p/|�B�=�c�X����O����X�'eBx��\ �����
Q��7(��ta2�\��{C�g!?���`{��&W!�j{C��� B���YSo��KOw�����[�x�o
�s����k�!�o��V� Ѕ���q��;����t�{���o��O�W� �1�+��a?TM��iL{������jB��n��pP�]�9�
B��UX�6�(
�����s��*�z=1��rWx��>�e�\��cQ��%��@��>8L��r���=����BHm+�F -�o+��܀LPɄ|�)��C̴��A!t4�r�n�,J!��:nV�#| �fR)Q�#�i�!:a&�]��%��0�gsͽ���*TU�D�ȹ�_Ai/�pR�M��=Q_]Sᕰ�x�[���i�9�!��<�!.���V���lb�Y�q`� [��߉�RB�c��ゕ_�7�B�V����UX�v��p/�� MVc#�),R��N�W��`L���`��kB�
�G[��B0,gR���T�b���ڄB�'�.⽠),l�+�.Z�����
��a#�O��܅p{�����i���&�L�B��@�m�6���p����\;6��1�7l�Bn$�{���K�k� *���y�y&�G�}���f���'���SS��Ы��P���`s`��r���.���so9��;�c�de����˩��A�r!�3�_��3�P��L�0�v�4� �#���t��?(v-=�p0���>��&��/��Jt	A�8Uu󔏣�>hz��P�н����@��J��{q}t]p�(��[���
.s�����+t��B�1���GK��2~��ޝ��p{�w�!���)���P!��|b��Nʜ�%�l�YA�'W��&�*愜H�B�����/�B��.��/,U)���I�@nX^�fa�H�rW���@t$�Z
A�$�����'*�J�&�\��݅�(��2�y���R�|��ҪD.�
�ݭB���و��%�s{TU
"�p��XMn⩒�h,'B>ȥ���dT�{G�1)�:��w��/�B������>�.(�a�@S�C#Z�Gter����B��t��x%�!�'e�Ю�x"�jԨ�@x����5���.���Bx"��FCɼ��;SV��op�*�}߰�A~5�,��{�A�޿P�N.ď��l���s��8��$䛌��3y�� ��������ˁ0�zCOt��D=:�����B�B�&,�>:����C8���Q��.U���C�.��+et�.񣡢���gᵡuB��U�*���#ر�| 8�5�~� ��B�uG�h��W�F����T~!�h������R�'xcPb��):�gB�|�j(�o!����w'c��!�	3࿪�q�"!ߑ�\Ȼp�k��7b"�\Sa��t0*K��T;'r ��³S��qN�ׄ#���9!��t_!�b{����,
a*L�M��z���L�Un��z7��
�*�e�X��O<п�؞�e"����d��W�a��`:V�]�GYB�M���[c�KME��Bx"5���BP��Y�s�B��`$�Xܰ���l��^�~�90��TR`�
����c�C��-��ڰ�	aDox��h5�D�|�K��m܋��wb!Lw!ܞ��F�n!v����M]noL�wu!,`; ��u�U�s6G�?@-��B�梃��B���ɫ��y�j��Z�r^��z��9�3~�ar��y��q�?BH�0L��B�b������Y��H;�O��� HN*�	h
'��>H61?$�Mp/*�O��G��C�7S��O��B�LAbP�i�
��A�ƄP������Pj4:��[,��@��rq#b辁B�>Bք��dDbn��`�Z�m/���%�7G�(�9;�D2&!Q�h�pb��KSR�υ��jzn,�����ى�;tt����"�!���`G#f0�EjTR	��q�9H#�����d>�O�� ��v��!R�Ty��;���@���ϴɬ}�ځ\���U��;z>���+^�٪ߌ�0&&$�|U�;"�����
��j6d8�b��o���_8�q	�n���*�_��5~�����_��h�r�7+�#h���Oa6~�EW����p�3Q2��f�9r����!�"
���1�{�$yٔ�DX�g��p��}cLt�w��"��؏�����E�z&�=�ّ|ov��rT ����Y���Y���p�Q>�ވ���Yc 7��1���
ѫ�JB���J's�Mm���3�)́M�����|�z!�c`1�B#���y2LC��0s@S��O+��I�Y���\�soE0���enb�4k�#����l�M&<6�|;/��:��Vv1��7xsRb΁�9�6'W�	{�f��1�Q�4k6�*�h���D��dƱ9y���ω��JІ{�oO竄�EX;&�̅s>!ȉ�!��E!��0O`�X�a�㽺��3�~�|[Ś?����x!�A�y����BӊNBG�j=�{j&��U�Bx��2!����܈����2zsLl��B��^������)�|!����B��{a	�HA47v�Bl��>�M��z$�� 6�y������,%i�NǓy�$�1V��n߰�=�/����p�����w��X��r#�|U����P�æ��A�0
���|Uù�I6	�
�;ri:T���|<���T�Zj�E
�x�eK�����K
�kbO Lv��qTZ9Mq/8i��5���S�e�(��	aD3��$SP2�/#$&�?	���HH�@�!#����^�\<Br��L%e+_;� ��"�*���W�TD*&�v"�Q�&�L/B�'�^*�=���B؊$�K��C+L"���Dv!hi�<�39;�����N"�G�MIN��&L"ϼ@b�xݹK@r'�p�(d�*Ϙ�!��Q��&�Z��ƾR>7G����m!_t���c�|"�����P�iSC��	����{@#?B��E�~/��ۅ��B>�\Ǭm-��G!6"}B�X𦐏��L	�!��j�I��ݘZO�Nz5ĺU��Ŝ]B|G�3Z���2qav4�6��Y���DX�+�n�r!4�Bn$r�W}��Bx"����C�>\�YG�A����3!_�V\�+WEbG�!�6a|u��,f����L�UHIQ�_�ñ��r{�b��ᚕ��b���Ս{�K�|Bѫ�j� � `��}��o�I[k^���B������0�pNb�|��v�k�lN�OM!��Z03m�<��+����1��d�rk ��ⱅ��Dz!�x���@���{�2���:#�UF��$Q���BX2'Lu��1IԚ�&tj���';'��O��B�����v,@��� V)M��\f�OT�7���]�k�X_*�B־�p��U�5����q���BнT�{�{�B���'ʋM�)�����a��J���S�X8���Ph*����JB�CL�Tȟ�a])��P�A�M)������gB~�-��aU�Ng�gKC����kS�m��}��0Y���O࢟�b����X�B M!tE����D�A	`!���0���*z��y��:(�T�{�i�4�1�J�	��l/����I��	>ڙ gb��K^�^Hj*ď����qO\|!T;�By�n��(�X�C���n� �\s�P<�{!oW��X�@��s�P��t�
�2�jI�[ ���]�2�מ�IR-
a��\A�1h�½��>A��Z\<�Y��!���WX悫{ ���?1QZ]��*���9i%K$![t���1��f%W�D��bʦŢ���B�I�%ī�z�
�W��LU#z�`��p7���P�B�h��H��MxP	�s����P&r�\J���HTO*d���ȅx�wt!�Е�J:���|��y� ��|��X���,�F��MT��|�T�A�n�B��m'��V�
��ۭdB>V7s*mV)��#jF�_��\��']�U�0b솈q!�0B�h+��B.s�>��n�-��A�evC$�f
��8�V�ʆ���>L!r�`05�
��8v�,ñYsc7�o7m�A�C��U!}_%|� s:��͒���;��)�:��7��v�B�I!�aS�O�U���b��H AlwxF������J��'"��f�!H�>��'�BG���J��_�}7]�+f-�_vG�q`�=��8�u�����*���rfA�w��i�o?�=˩T�\�0�����>�a�nA���=�{P������,��H#��!|ǁ�,!��a�����#UM�+��s���I�-�{�a��h���]����"=gb�'��8cP�{b��ٞ(z'��8��+�
J�D ��H�#a5ᗶ'��6Vv�La|1Q���D\f!��L���Wa�M��A	\�6��E��pظ
�
�*�B�,$u� ���T�rN/{!]�6"n�/�{!�H���_�kqw���-l�x{���X�JWIvЅr>{Q-����L!�څ�d�Y����\�_ |퍤̛gM{#�I!��{#�t?��&�Yw~�'"���MBa#��ވ��;"����yS�b܉:��`�$恇�f}�zE�� L!,`�����yp{��RGsxm��<�����4K�G3��օ� �v�(<p��	����b2&!?}(�wD�%�KȜ��Ap�f��>(,ā�3!���Z 0L��W�3uG�B���B�A�+\UG�> )�
��.a��-hg�	I�wwB��A��uE
�W)Wc�'p�#e>h�$���B �	�驐�5	q ��0��\݃�vpC�1��`�LD�	a�%`���+&��wNv(�8|!��\/��R�ڨ�%��aN��s�k'�����M���B�T�scMKo$�T���t6K�a�UXE��������a����@.� _���]�U>
χ�X�w<<��\����� )i�mbO��Cȇ�y�X}{��B7�
�E���)�x��B�!��� ?<E���aQ���Da	��.�}ߠ)�R#���o��wN�m��=�;X���T$�>�6OCM!�5]�L#J���z��x/~���څ||�GY�φ��B�&z��,S[+�'�>����@xm��:UQ/ԑ<��wa�?�FaǺ}:���"-�^��}����
a�w�1OG���b�D�	��
�B�����1O!��4�wݷ���W�k7�
�h�d��b�B����(^I����aLD
��(�v�3�z�̟��=g���8�/�]ȓ!��:���z�ޝg�Bh�'an����e�A�P��0�ک��@~
^F�#���ܦP/׾�tlB
<X*��m!��@�NXa�DV"!�Ve�+�� �:§��;ч�R>>rX�^�kRi�(Aw&jy��8̪v*U�#�ׄ�'��Z�{!z@ȭ��r� a�3�Z!�	n�܊!	0�����ވ�*݅��:��jn.:,k�T��
ۇ5��ѱ����//�81���½(��_��̗Bn�>L�V�o��`���h��FR����`Y��x���ㅐ��j��Ȭz6ux�%�w?n{r�b!o�F���4qgs*l*�'�BLag#�0ְb��L���M�g#y�����>m��hd�*h�A�g�v���V��X�0�U>3�_φ��lı
A��'�l�9p$(�/t�(��k��b�|h%;���:L9W��x/|ڃd���|ul��$O��8p�*�{-~��<	��A2�B�=*��UrIC���υ����'`9�������-!����N'(��8��z|�@*!@�֕��N��ҼƳ�üw�%PN�Ӳމ�	τ���L����mMv���!��DU`!6q��O�i3��%�{��;In2Is��$�L�v�@�'���!������BP�	[N"?�V�L_X�C���u 
B>|�|�I&�>��.�=!�u!�� =�D�/�� !v���!W�I����J��_��M�%��+B�r!*I�)!��B��q�S���k�BS�$J���'�80�"�s;V�BWyO4�F�W��8a�)�*�
bS�s*��VL�v�K���Ѱ
񅠸	a6�j���OӪA��(lpC�v '��`�!��GKw�r=Z��!!�#ܥ�#h":"$�U��^p��x�����\�fQ_�#�^!m�xℌ���r�����Bh=B�˱�W�]8E�w.���5:JAA���͂7B�$���F�#�zuPb�)r��f�9R*9F�@i�\�Ro�k ���ŽPGS��ׄ>�O;PIȵ�Bh=�c ڢ�?�����.*��sE�ڋ���,�zL���;����k�14��H3��7��N��	��@!^��
��|��xw!�"�D�v!w!����b��:�^�Ф\�0�Ą�\�i�*&�R���O��K�d��R���R��'���91Q� �OOkb��Y�]Ղ��b�y)Xʦ�B!t��Q|U{�O�֎�rcB�iJ*�����RΒ�B�:r�A,�����d}w!��c�D-�Fpo�]��k�a�m��bÑ����G���w��
���|܄���bsLl���e!�cb��+i���	�r���<y� s6��	a�gb:!lE�g���8p����!rl��7����u;8)���Iyq8��V0\!<q�'��1��x�-��9�X�z$xG��ȇj'��� Ig!�i���98��|<	P� ~G�DyS�� �B"Ԩ�	^0�����U���Dx�+��^�(\2DX;����z"(%��s��"p�U�pj�)p��	G�*̓�t.�����$B�/!�}"AW�V��
�\�:@"�RU��J���,$��À"Q�L�/�YX�
~"�N��D�F}F�6*�U��©�i�	a�%7�X7!�Z��H�`B^!����+�w�1��0��\ K5�����V�	��j&�5]�5�/��&!�B~Wu��z�rQ��K��	�*�$��Bh
!
�'����ɓ�d���ᆐ�{)�.�ܨ$�.l�.%�+_!���6R����{x�ū��	��7RB|m�,��5BnȆ-e2'��#䲰���l�x
�drM�Z��]Z�0
;6,��qB�d&Cw�ЮN�֛��p��w����Z�P���ʊ4�3�r�@�"Gv2�G�u9!ю�vvy's�	a`
�s�f#���KY�u�_�e�[x!��!~G�WJ?�t�Pa�/C�VQ�qr�Z��@�9!�׀����hng���ޮ��K!��;y!� iJ��A�b���{��v]�'3�%���0|\�
�ȅ(�G�`�Pa��B��,mh 3N�P�z�Q�Q���-!����s惩0����5�I�ٕ� �h��M�+�{�Z�~pW�d�!!�i�i�NM�[��	Cw�0&&��D�UB?,��d͠d͠�|'ׅ��i���d
����<�Ʌ��ʷ��P:��BDoyB�`ͅƹ�Y5�mf�˅JB�rl��7���(5���Y\�(F��%������\\���B�!L�����^v����v�g�B�����F�!|���B����k#�P��F`nnT�(�'��kb.H�k��#��B��t���p#�o�LG+�撹)7�
�%�����:8�΃B�B��^�B��<2��cDR½�5Ы�����xG�P
������C�ơx`�σ�y(W�rN��N� ��?���:\�`��<��Go(��G��w:� D���� t��,�j@Hq�,�S�@J�B>�����F��$;�Ha�s�B�=��Tyw��-&�+k7�B��S �@X��=ydT?D�R!l�)��C���_��ݒq:���B����(�� *lR9Mԯ�D�L���q�.Q��L��D<_!ܞ�D*�B�B����$i�Oxa�+�H�!Q��r��^8�/����xT���.�dh���kZ^����7j��� ���/��X�� ��M������.�J���|�[;�q����ܛb���|�Yq��x�;�ߌm���m���x�kx��7�ny��oy�ɋ}���_�c��t�/6?������=���b��-��q=�/ˏ�݌�/�n���{��bmi����Ǹo� ��>�K|��?�w+�\v�����o�����79�����ƾ��/F��n2�K��S/ƹ�Ng[�G��|�~͡/����'�6x�k?x��~��_����G�'�e_�-�}Q��͹����n��~8�_uz.��9/���_��˒�\�ۗ��=����i��U/�����N��u$�b���s���o9:�y�T�/�q?�o�ew��b��19NǭH�b\S��:8&���8������196u�qkN������� ��Ǹg��`����8�_gC/��������b���&�~3��|�1��oo��Q��,���w�7��m��s��q���{~��f�|3>wrl�ɱ�:k�lQϞ�ccn��Wz��07����ҋQ����<�Y_��^����yR��W�5t�G_��c<�o̤�Z�}�>��\�נ>�
�y��g�k�����������ӎ�&�㰽�H��Bd��ί���AҲ����{�&��c~���+�k�W>ק�6)o�������|޲;�+o��U�^?�z��o���k���k�?_w�{��f��s�'�����z������p�/n6�a�i��p������m�I��R_���c�و_o�5���X�>�-	�!���u8��s%�^�������yA^=K����X��9>��N����m^K�}�#�-�>?����}5�u��!��5?f�\�S�U�����s<|йѫ�n��{���R��=��I��C^�[���N]�!C���9�l�1��c��O�ۊ�v�9����k��f�W;��s<�S[��������Vc����Z���>z��^B >����UI�- ��<�㻟��zzΏ�_σ�=p������W�|��-���c}�χΰ��J��2f�ն��La���jҞ����m���|M}���s�|^�ro�W.vHU��L~U�}5>5�?��N�������=8������B�Ĺ8�[��Q���1;�CX��0�&��i�p��}h#�u���9:W����§=?ǫT�nڪ��iAA��G�߿����������������Ϯ����������Ͼ�����T�����M�?�S ��7�nE�?�O��@��[��On*����O����k���:�:=�ǯ��H���K���4�#��#�U��ߦ�ܮ��忺��?��Y�ם�< ��haN��_Y~�q2Ӊ߹_��G��ꦋ��m=�����~�C�H���{�x��p�7��������c�ߓ�A��^�z#W8	�ո��{���H����ڏx��d������Y7��%~��^�#x��!�Ȳ>|Y���u����Ƴ\⿊n홏�ؼ;���2�q��a_yެ�?2'�fʜ>��ͺ�G�?�Zz~dO'x�M�#��9>�M��#aw^���z�Ϋm���.�V_d:񱺆��>^V�Y����b-_����w񱺶�U-����}��>/^�u~�{ϧ��u���!��?�icM��e�n>~v��a�Д?���v�o�����M��5n� �I\�:��J��@�G�~O��H�J�����w�g��V;Ы�wC�ع�7��Kj���]�kϹF��7}���	�&�������+�+5Ώ�t�~�K�3]oy%��_�r��@�|���#=�~6���8|U�ğ~���:Ɂl��˟�h�=����2���hN\�Fs�;��h����j��?�v� 1|}�{��G���W*�qi�W�Xއ�|7�W�W��?��� Z.{#𦷎Ώ�L��yZ�<����� ���l��esM&!mR��]��hI��	�w�>ss�V��eBNϹ�[�B�a�I����Tğ�}��5�G�{�<hO��ח�G\>g����@��m@�������.�w������uM�Sq��x�ܩ�Z����A�Q!b�.��De�CS(&䱜�Aڏ� ��I����^�y:�ƴ2�i�ۃ��B�P�b���<7DcZ��E�"�	VK��؞�P�[c�!RPȣPZC$����>B�.�ʺ
a�6j�B�D�'Y�<U)��#4S����P�����c"���ۑ���<?/BG�>k;�5��<�M��ڞKC��Ʉ<�:u`��T)q�6"�+�
��-!���q{m4Cj���*�`�('!�10��v�y M]艁[�D��$�Ib##�=B��D�m �j�����c�KĶ��}��'����y�;N��X�p/$�mA�����X�U�������Z!���'h�VBW%�1)}'����l���X�0�gz��BhRY��W-T�-�M]ȟX�G�<!�;�(�
e����B��ƒ�B���@2-$.�R�O�Pм-������oט�Η����m��h��Y�_{�����mOl �1�BX6Rc6f�.�{�lJ��c�0��A#z/э��B�����]j�>��Q��l��m̾]�B`�D(�y������O��|�-���*z:>�AZ�v��pou��CK�T_��R:� L�ʻ@�/Ģ��e�P�:ǃ�ۡ:�B/E�$�С�9��C�>=���v<�'��
d��>�ه�x/�)�q���*��y9
�]��@�y!(n���-?.�'"#h�&A�TO\���H-�vM�I eg�$ݎ��ʑ�UIi�ȯ"U1��1��%��� �i,
yO���B�W�Zr�B4Q�Ei�։t$BPNyrz9C9j>�*wi��П�O���j�@>a
���?ZP�?�[��t!�������˿�2��Ul*R�
�n����4c�%����R������UQ�5��j�������� �L���je��QC�w�E����	zC���B��B�Wx�$!�jx�[�U.s�\9�!�}�Q����?��0�:R����W+uH�{N%!���Bn&-��)ӭ\���[�j%�j��K?����/��Cqr��K��b���L�c��xeh��(v$YH+Yg��B���M!W� r�Iu�;�J����{������E��;��E�cگ�\���x#��1�\ȷ���3!�D5�1&�p�]��9�'�U���*��CH߉���/ĥ|���d��!U��y��D�r!���}=���AI_HWb}�.��	��;���YSt��^���zl݄0�6�R����A�P�<v�����zuA�.����o�;���u�Q�O�=q0���A�-ʯ����7L���s�u��H!���ߴb�H\��~O"2�Z��=Mk4��.�Q�^ru#KY���o.:��B�/�+� �����B����v� :��2��v�p��[��g�V��}&F�~�ܻB|!��+w�·�A�δ�Br���x{���@��B��hhD4��@��Bx"\cz��a%�^���H������ �)5څ��=��$&�̖Y����| 1�օp�DU��Dƽ`��ܻ=Q籐Gڿ
�GKP�Lg)�&QͶ^�{���hR�q��)Z�|�l�'N���Z�|TV=GpJ�O�]S!���x��J�'�w�v�ll�T�p/�Ǫ���ùdЖ&�F���驐�4!�0�_(\�b�����f�����hH^9@��I�G�1���@�
��b��va[3hgt�-ш�c��J��C�x������ۃ!�}G�Ma��&����&���c!��|BLʼ�}-�P̡���()���	���9��6Q!W1ƀ;�X�� �� ���*Y�v�|��B݉1q�$��)u�o?��֕g��l��Ӈʰ��vr"�����j�[j��^'ҫ0L�@!ܞ6!|��ܤ/������C�r�U/����I��/�p43\Z�*>�K�
���Ocs`�*�F����nn�(�B�p���H�O��PɄ0;6|܄��ǛB�c��:��U���|܋��������C��{�')��u�1XdH�'��F���}`�BOp�[�_��J�:破��ټ�6�eƁe~���^�Ѩ�9.N�%�G�xsջ�_��*Z�����*��3U�h�D�96t����`�pv�V#ҭ�BlD���S(ge�| ���#'fmR-Ȏ���V�N�>�p��{������*M�WsC<j[����P�2'�u$��-T�Ck��4ѕ�v��n>�:��;��oh>ͿP���Q�� BSQR�P y����h�� ���Q!^�I�=��|p�)�S�'�l8���B���6]P�|U���_U�f������f�~�+x5�ׄ�nR)�}�7ؿ�\bζ�9ۗ�B�����L{4�l�n�W���fm��]�g-��}v��&�K&�:�00;$�^����@��a8��?�>���~
� ��FKm2!z�vr�w��́�Ms���1P�L�F��	�,cF�@�X!|�1\%Ӧ#G[|�~Bb��c�9&+��U����7��W�T�r� �6��!7vU�t^)��ÿ#���\�%����(�Xَ�ClO'#���_6�9q|.�V!�Չ��sf�WӅ�'���y�>���5���nK�w\PN�|w"Ed����w\��
A<.�ǅ"�������F`S՟����ڱ4!�O���0YͶ�7u?��踊�ܦ�q�S�Gؔ֡�!j�,Q������|�FO<����J>�{�^��ڃ�B��C����^	Ӽ�g�ɢ�7�`�)e��?S!����ِ�gcp�i�Fߟ�tp�'����5F��{�uW���
рA* ��h��⽺�U^��3`����,�ps�1�3���U��^ܱBn˅ME��v�q�.EϤ��~�]��h�d �QFB��90�rBJ�����3_9y.¬e��L�|L�e.q�V'F�p�|Z����j�
L��p]����~�|D�i7}�G!�����"��B8�XZq�=|��a�<-W�w���cU� 4U��;��fU�ø
���`�\5\W��N%�;�豐�|��T�#WKv!�ri�'��1��&�jT9>㇈b�kw�}�|a]���mB.営�hD`Ltl)WGނ���ks�v��
�dZ~V�¯pC-�=1�H���v�7!��1\���*��"t1����ۣ�8�r)�@����W�[\���B_�j��횈�BQ�'G���B�۵�v�pg!׶�,�|�!�Egn�5�W����]�__���i'�����ڵ���ֱ��B�V����v��څ��EW����v�o)�>$�
�R�q�)Aĕӵ�-��a`��1��n �揵8 V��C���G�1B��_�v��a
.�M�p	�N�v��]��m���@��JJ*٦ڹ�7jm8�Wn^��b�!橑:��PO�w?��6
+�N��p@�?�������JG�'R=�`{*��`oU�_h|�0i�Xg�n1�K�v4�`����$& �?�I̡ψ~���9[#��8)+�wtP�	D�a�	��%0�_�1
Gl�iBx!x�U�,�+��rZ��\M伩�_@p��>��6}�r�%P
��Cx�a�rN�	ÄS�����������k?ر��8 ������~�kS�+������/F-|hF�>�>|n:H��٥o�#gӥB��K��|�B��]B>|�^H�TȻ��-���'.�U,��^�7RB.�6}1vC�ޮ�s������\��vL=υ{�Ģ'�סBh*�B�b��`�t��x/����2�C�،���c��;:w����.��q�/�.�𪓊��c!����c>���Bl��n�M���j!�r��k�D��rmHȵ!i�lׄ���;�+H�<��eV�8~���*�{A%��B��m&�r5j3CnՉ�F��)�v�<lo�|�U?��(�:S!4uA��VDL�Z�&�=�*��^�B��T?�����B"���B�|�H�Q�Q����{Q�黨�,(�BnAڋfA��̐���M���AU1&ޅ��S/�{5wJ�8�S�`�m�*�4����k1����]v��C~Ǎx��8��ὶ7�X+&�k��8��������F.�BhjB�0�
A(��7RB�0��w<�r��f
ۊN��>�:*!z8LR����}��fӰ!�T��&Z�{�&�B�!�P�0L�v����m&�B�c��Z�`��5Ʊ>2�Ď��<;�U ��D�m�*����pKڌ��Z��[�4H��%��o��H ������$��e��8Wª�TD1B��0/�{�N����ba�����f�\Ar�>ã7+�7:'�GN��DT��߫�7����@��9W!��<�Uz��h���p�#�_!����΃t3B.:�܊�5�儐�m!��J!s� �n!��aB��0�B�r+�[����.���ą�B�RN��!�o�۷Ǘ9!�D��?m�(�M%��s-���`hhX݅0L�&!��p��ƿvC$�i����*�#��a	'!�s�0V;�	�V���vG���Hx:��-H�ՓA���hRa��t�
!��G�U!4uP<o��1��P�E_h���T: ׬��b���h!|G�Ԝ�g HN�7,B�=�q�|Z�w�w����CO!L��Y3��x΄��H�]�3�D���_{��^�"B�(|��jhS��X�* ��8�<yϢ$_]�=�^��Q�B��YH�qV@�X�_���C��a�m�ர �B���m�	�ko�=1�7�ꦲ��G>{����$aӦOD�Tm�1��9Ay�}�Tu:y�j��?�F#� �W��X�BxGΎ��TՕ�UV����=�lF�F�A%;��'��3�Dk;��-5:f�鸐�P �� ��B�ws�x"ұU�^妧�*w}�[������Nb�&394�a�ه�B�W�HH9V����V�B�tro�Юı�a�ѓ0�i�b0%j���kv�c��K��+�^S!���$��*����I�S�n���{�[�Llu3}���U�~9BZP!�_���]��!���p{dLr�[ɒ�C�<���n�l�B���$�)�����U�������Ѧ�
�T����%��B��\�����[�h�r���A璨rf@.�
�lj�RS�����ܾÝ��l���v�m$:�{!�
�!�r4�\��6G�oz�̋�}�'��<T��V�q����-=���x�ЅLRȇ�@	��矶���N'R$W�,~8\rmHZ���1��B�W�?�T?B���# s
�ŀI�����5�)�ؘ�/��a L8��D"�J���8q<�p��zx!d���H�$ĞXn�	���p`���~B�$$��:����d��a�D;&��Aʱ"M%&�@���؂K����cQ,�bHG��P�X�kQAZ�fA�p�^]H�QM�g},���������oH���Xp{��ˎ����\N6�	a�l��Ħ�$+�1OD%!���}+���k�4�����d�F���IL�f�&1Bl*����cՄ���Ashsc�)�6ibs�۰�a��8,�}ϰ�8��
�2ڕy�q��8K���Y*�x/jCu���p�s��ae�`�U�&���.;)�.q��9������@�0ږ{#�~"ڋ�Y�Z(��l��@E��*�}8b�@�:-n/�
�����U�BA�4I�M�ZK'!(H��G��d���j�M{��Pɘ5Fc"�Wu����*l"��[����1!���`!v4��a 0)M��m�䶎d��B仦B�
�s!�CB>E�|��qB>|�'p4#�ӽ~$M!�>T�$���
�^�ZQ�W���j�*�]H�^9��]�&K�H&�F�~��r����H��NfΆ�`!�jìM:	%k	�4I&򵣤#���\�����^���V2>��(��;6B�W�k��U�6$�ƈ�(�"���Q�E#�#
W���;^vxY��Qg.�9z��#�+X��״d=i!?�́#�B��{!<q��*���Ѕ>nI�Yx���.�t("B� ��IMMW;��1Q�[���9���M�u)�`"�h2�K��VI[ZV�^G�Ή���ۣ�P!��ʫv!���(%�Z�V��㔜ȼ$�):�.��w�B�Bޮ��KB���p����\��±�4E7ޔ����(���'Y��Z��
��D���Q�Q�B��i���[����ڍ�2��8I��&2��ZB�]$�vw,:t��G�0�V�����dȚ��IsS�o�4A2m�
%��N
���q�-��}#L��*���B�w�m���@�H�QM�џ $�A ����½p$�}�l/%� �uҲ��F	A~�3≨9�!Z����[$��ɃC�du�,w v��GK�+A���$i����BXQYB��GNԵ��~(������ض3�O�P&��
�*��@�d<�&�]B�>$�݅0��2aCN��U�����$���93�#�,�O�J�u(Qt����p
-�^;���[�?���T��//��+�^�f\v�o6�nP�e�w_l�7n���ȸ얩}�_����`���o��X�`l_��܋����W�f�{��q��3��}��v�&_l���-k�b��6:�Fm�V�;��Wʣ[|��x�=���J�K>#�4�/����L�	�^l�{�'�n��[�+c_�����b�֯W�eW׾l��dr����s��d\���30������3�s�'eNϏ>M����^l���x~��~��w��}�s�����b�c�c��㺏���X�?��f�x1ʿW�������_l�=�su��~N��q���|����Ÿ��~���b\���:8'�<��oo}����(O�f?�M�87��ys|��w8N_)�_�c��p�|�\_��.ˏo��3?�GR��d[�����r�eV{3ޯQF�ƹ���j��v������[�~�f�߭|�b�-���ua�_����������2���.��p?إ����,���	��!�����7u^M�I��/�ۤ�_���ݽ҅s�d�������W�{�v�n�ͅ��6~ޯ����P|P�j~����bm������ʸ�K_p����߮[�߽K\�Ay�N����ԥxz�V��=7_3n���r=����������<�?o7��5B����2ۼz�����_�����Z�?�º�������=����+����=��r��>�m�=����Q�n�諓Gr�%�6)nʵ�𾙦^]�85�;�|�C�	��<�_��:��:�������LŸn��Q�x�X�"oM�וχX{�r|͎�N/C���Aݮ�������c����{0ʐW�z��87���|�G7[��_����ٟ=�һ�ʸ��ǻ��p�����s|���#M��as%�z������!����������������ߪ���OQ�\�����~r�����a��O�~���?�{��͟������.���%�a�q]=~�:�n�����^��h֎����.y������/��\�d9�����d;���?2��O����vP?�N�j.��n����t�?k�Mo��Y���R�#��|dzo�Qp��9�?7[�x?�\�~d'�;�d;��)?��*3�#��p��߫_��K���g}�W��q=n�ȭ��#�w�H��揜��\w�?�O�W��os���s�U!�G��x�{��[��[����`����=6n~�?���_��~$lƽbY���n^�?2�^�,�Y�����#���#��}������?�2a�JW��?�����w����ޝ�����ڍ�H��5���ٶ?�F������]�͛���y��r~ސ�?r����>N|h��k�˱y������{��.�k�ϔy\>W�j'.�����8��sybmZ��z��{=~�uc��5��\sX�IV�q����.��(�_���Uf-�U=ω���}�V].#���e��ۓ��t�����4\�\f�_A��� �����G�+��i/�{��ڷ4�%��{o������K�}��~����6��M��d��O�*w��9���yV:�p���WݺKH8�oz0+Oǳ:�ܽ�^Nl�Fg��hN����9x0���=�+��@��G�5�3�De8t�#�,_��v�v����8����%�ԯ	|�pis#*ph�'}���Wh��j�y��W~�k�#���G|��XL�y�l��N|d�����M�s�?r|ԉ�}���>�"\�E���t]"�#}l֝Hu��c��n+��y=
~�W�쮽gw���w@�p��ܮG%z>�G%�z�$
�w�0|�e�z��3%�����?�%�#3��Gī�I��ۚ��>��r�h�r�!���9����
 �v�!���|�ۂ��� :�n�u�O�{!���'�r����_�=�ۃ��B���'�s{�MW�_�/�8�?Z{<%�zU�?mCݶ֐�Dc�u���iS�]ODa"!|톜6ux�{!�`k���y���o�C�j9��i[z~	!�/������蛹㴐�(yT�z�#dH��9L�#O�����Vy�GfhĹ{��GJi����Б�³�C̴��g!��1�0�;R����b��!��#pM�-�A�1��@�p4w��6�i�
a�Dy����B����B�
E/� �Ɔ��քw<X�*pց��*��wBO �o(�Q���Cf��j�z B�91=B�:XH@f"1�����B��&*�
y�`���^HV"�):!�&WmyѮ�^��`�!�jbS9 &�#a�-�z��k�E�b{q�.$g⽐�L]���Z����º6$�B��PNJ���)�11�� Æ�ڵ�|���aLld����ֿ�7uw>���FNT!H��}���3�Fn"!Lf���i�{y�_!�{���AR�p�������F��Bh*��½PGQ��@�BxG��ma�BWaMcƺv���	�Jմӱ"��lg@�>�j���!�`�9H�X���!�ą�C.�@Fn��"!���(��i���)�����R�[H��*�8��lHBX��Z[����j� �Dj��Ņp�	KMp�2�����f�7������w*GD���������C.�^��J�p���D#���H�(䟶�rA�g�.�(�\���C�R��);d!K���b(y��F��Bx��0���%�4Q��UJG�U��LZr���2���՟�eN`�r�?P�
5 A�\<�g���4m
�	��BٟŦ.���}�)���S��˅h���;k~�#n���%;��(�i&��؟��W(����X�W����a���YB���y��u�&�ªӘ�_��?��W�A.�ݰ��rB}�`�/���Mo���!�պ7$pr5�����'zC���*��C_��j��\�
��w��娅\U�e؅ ��ժ��D�0�&E�"���+�1�7&_G�!O�i&�]+WQ(t�B¬�Yؑ�^S��2/䆠2Z��ҭ	�Y�7���gm�B����$C�i ?t���;d�z��5�S�\��R��ą�#��#���	�
�H�#�Z����@ٛ�
X�ȭ+�x/W���i`��tz��^���g�{b"�:g"�u�o�쐘�>a���V�څ�(�x�o)��_/��:�3�,��'zV�V<�;�0Eg�]��('�+?�X( �Ut5��B��.�Կ�����GK�E�(s�}�(�����0���_{M����B�^}!���Jv4��B� �`?�N�o���ºQV�w���;V!�
�W7�\�+��B|G���#\�ɵK��kSl��	am���>(����Ы�!��B�
fR!��U ;+�V|ncD!�6R�	A(����qPհTL�*�靕z�I�'�\T���O.�g�΂�=��ʰw@;S)
aw��^&��ʅ����(��S/J�X�	�qI�����v�5Hj�@�e.�*��\��dN�l}g�!6"�B����5�3-�YϤ���O�i,�_(q�#y���Պ��Hdt�4�
a���U!��Pzr�(+���[��Z�O������+d]8X�DȕS!�B>�j�� ��Τ+kH:�.'ƃ���A��*-��|Qey�U(^"��x��{!�rB�9�s��0h9�hR���Y9�z�2.FC��2<���q�����k
����K��+���B�<aȱ\J�⇰�W�X��W�Ѡ�W���h�0 ��
a|58��WX�ai*�{!��h�����{m�.�hІ�+3�EW����ul2���_��)'�:::EG���
��8:]��Ѵ�
aZu��A�v��$���({�gsB�n��D�c�=��#�k��~ �a��ڣ^h@��=���(�@!:!_X�|E� ��H-��>��� �^��.bO �o х0�^a��'P|I����B�|��+�T�loĄӱV���_!���B���p5��&p
yM�5z!�&�y
�*H�	k��'x�.�cn���B�i!�W��� �&G���ȬqS�
>�X�f,*5�c�[��U9s}���f��h�B9�t[�D�7�#��,�	�����z����`]�h��܋`�8Es���B|"��4A�7<Im��x��!�7|ܴt��5�$W-?�*�FPǤ��x�_�%@S�BTC!�BtC�xܨ�96��_���/�ޤU�?D�*!L��v�Ѹl�B�گ����9%��3�o����
xߑ���	�&'���
s���3ΠMT�6���Lu\뭏�{u�k�\�	��JeB�c`�
~ǠrJwϊ�iy���
x���*pv2ѮBX���@��A��3�>�&�(�*�,h�H���n������O:�}�n�Q��ÿ/��91�4���sA]I�	��`!�K�Hnk�#�V>	�h��b#�� �-%�I��g���u� *�Yȿ�|WY��D�ok��_!�',B>0烠���@�|��{!�:*{t�4C�Q�[��
��u�gE��Ӿ*�\�'6����ʄ�^8���p�P�B������C��ELgۮl	�J&�:�l�u��)L��|_��6;*�����"
���BO}�5�@b�3;�uTUoD\s����TB���R�c	�m0&^Y=/�T����À0;�'�B+��WANt��������D=;EGv!��'M��Ы؊́30!H���96U�Cx��}}�;���9`ȞF�*?C�+s,?���c�j�8��d��P=�(�V���'��=Qw��Q�uߊ4�U����:<'�(&�BX�'?��B���_�A���B��4
an��g:Bn.�=���D��qP��Йh/���\0+A�X�oԫ���:�_h5�m�P΅��B���XX�`��=�|�����R���N[Q�BŎ�*y�^A�O<�1+�n��r.�RV} �2��	9���I"��G!,`��B
���V���F	ֹ���I�Ua�B�K��
�_��-Ħ"�L�M���d}�&�hlO'����`<w@bn8 VA4t�K[σ�2!��1BM�B���Cbd�(�'v�|��r{�����/t�Ln�^	a�q�ǳ '�::\*�0�ρ:|(��k���hӄ���NBy8	)��蘵�y�n�U]�y�;��R�Bl����9R&�!�G3U;��w�t��0E���O��ٰ�$�����W!]֤����U��&L�BX��y*zb��j.�!��@zV��HD��<Xt�<B����˙��r��L(�A
�E�B�6�B�'_%��|M[��G�����`G���(�t'�B	�{�X��ä�O+!�6�TTj}\�tlB�v���B��UMO�W�Ơ2�{5H�B�2�
���p��j����&:��K_���)�BX�jX�0��bmW1V�QI�7׫��$�~NESå�6s�B�VU��(��Յ��a�t�ѯ��Ű���C��K���Co��i��Qq�@���#nN�u���D�s��п
�������B�a�*�Κ�|�[���|aC�נ���*ī ��i��� �u9!L�d&�����q�|��<f�]ۭ�k,�9#V9* �'�'�f!v4�#�ʱ�~>�.��\u8G�#g"xMج
�Savw]L�)�5�y;ל�rL�)���P(�|?T���h�f�ZPO��@rb7��n�Y$!t�47���>��֬�ve�Ľ��B�Ūq���&D�{xm&�\IC�/�?�B�<!���"n�̪���Bn��L�����h�F6T!|�Mm{��ƦLȍ��.t�I1���O�+�b~L!?Z^]!l~h^�8y�*��׆'ɢŭlϸ}b����p�t�4F@�π@>�:����r�0�u����|��_LM�N`�q
�A��bJ!�jP�
�h����B�B��M�n�Bn���4�MI!�GF@���x
����/�'n���8!��o�X�0�����Ɓ��>ȉ|��SWq�K8�a�&��+�E���-�{�k'B��;j�̞@��*xǫ�3��v�<X�`�0�J$���Q�\��L��W��@9r�q9��#|��8�x�/����)�-�M�\C��~�#��M+����BxGl����JO�B��B	į�BP܄8�Rȯ����O�ݐ)t�M����!
d�����~��
�!_ǦAO��n@��B>ݵ�@.'v�a�z��Q˛Y!7�B�����#���~��[�����t
��9�;<�����u��~�7m;|��Qr��(C�w�g��#*�	��!�����-!�	�����{��_�w�Bxǁ��!�B����/��
aD��N�Ϥ�Ѕ�n���\r+���[��;��½8 �6�@�+mk!'&��0�&�(syGOx�B#pޱi�r۶:z�ܭ�;�k"�C!�^uB���`�L��~�{"gj!4G {"�KZǢx\��	��#�Y�ЅQ�B��E
�k/��i����!��!��B�߽(P�k!T@�|�/��Rq��
B���!vl
e�½�0ood����qR�7ܥ6]���n��l�x{
��J {�DE%9D�0�7웕r��dn��a �i��*�]��%*��7��e
�w<p�ݧAԛ��>��hg f��#� �Wyz���x���������J�� ;��t7���
��A�f��ԙI҅�u�z�1 s�QBV�]S jF �K�.W�]����$�]=v�'PjAp��0ٝ�C��ODn��ɭn�Qe�{�l��=�Iw�e��I!�~i�EODĒT�DQ���ٝ���/M�=a&�tB�v�0 d`|e`�OW�B�9�AVH!�UI/� �Y�$�}�
�Jvh8��w�Q���Sȝ��\��{+!�σ�P�9>k�D!��J��B��B���
�a8;��"��6�.�NC~��� �a!9�����ߑ��MbB��4K�
���CǱCǱ����%v�*����s�U�! ����<[!>��#Y�a���R�B�VU��{��ڧ�.jOG���9�:l
��/����B���**����
����5n܀p��@CH��StpD�0��
Cn$d���J�O�:�U�����Պs�	�R^�1q�&;	�s&l�B�%S����p��LD�a�\�&����<,�q&W�	/mD\����7xBn�:�K�L74B��Vk�D��B�C���.C���)Ot х:R���UZ�{b�m�nO�$�'�2�a�ÌvBC&��$wg�!��&��7g��A���|5.�B1w!��7A!׶3�f�;�-�J�u���g#L3m#����F$��&�����Z?�$v6�����=º�)7�N
�^P}�C�|����qc;��V��zg#�I!�+�Y�b�9����R��}ځg�:�b�98()+l�B�,�|J8�j
���Q � ��	��$m��-Y�!a�
�oa�?Z 0��§e1d-���wX�̱v`A�$��TKy 9m�ע�0�T�/�*���5$��H�(��*�� ��|P]Ij�IE$�yX�X��Df	!�j"��I�>A�'�;CH��B�����u�ЅH�-��(9�*bG#%���)���N?s�G��|B��	��%������9!W��A�!7h��2Z�M��&B*���xW^��
��~���:�@���1��O[?ĆXȇ\мV�_�A	�% <\�\�
��E�UM�����*������*�EZ�r4�	�1��mc6���W8z���0�������P�^ȍp���ȍ4!
�B!�����Z0]��{u��]@y�{Oth�u��]���ţ�i��ͽ�!\w}�ћu��hP�җ,�YEּ��JB���HB&�+L0s��;��@<�>���1p���B�	��B#-&�*Fթ�!^!"]b`�F�
aZ���bP�d��Ό'Nd���a��q�p���U�ϻp"~H`±Gs{"�4~�2��6��Nx�Ąx�A#�����#|L�w��drBnp�������K���XpJ(��8&����X&���loڦa�p1G���	a�/D�Bl`Ж̪V�G���)e�����Fl`����6��cS��8����b!(H���B�[�B���W��DO�o������i�gqP�4�f���"^�'�b�q��J�}��Auz�{Й��Q&7"��_q(jBw���;p.�C��:}�ʭ�n�!H�@n��s�dA�WHr��-�}/��=ܝ��CH
��TW��,��0&~7ɫ�DB~?Zp�F��+�	-�	-��6��B��DE�B�B��!��D�?�5�c��Ie+��]kG�t�n��~!�ZVt��׆÷��ބ0�i%���S��7Ï��0�X�V��J�C	�E!������45��B�l�sd�6%�p{*�'�2{*�2G��|P6N�媐�ڤ-M;d��%s�	�z'ľG�������\���]f2^4��$k�
�����ޫ�g�x�l��LB��TH\��9!W(����K���Ӎ�%C��tsw!4Un�]pKJ��4�}��U���x"�M�x8^���p�t\�{�B��	a`��"KEv��r�4�	�Y�킃��eN
?��#����]7�D�XJ�����ˉFNG|2hU�5�Bh*�t�c�%�ۑ;2ihB#��!B��BYW!"Ns{t�ꀓ�>����n�)�F����gxV�N ?�HƱ怕?Y�؀0|'�?Ձ��~�KL��C�r �&�&�OT�^���Js8B���$����i��פ�����Bh<6r"�^N���a6i�KZ�
}\��U�n��s�����R��Ǘ���Ȼp����
X��{��Z8���P�֠0Gj'�i��VJ�B�z.
��Z�2���x*�WQ�X����E#Z���aiN�}(�#g?x�FA��k_n�/-�v7�G��~Oэ��B|���X6b����Q�bi2�T�� �b!���<�O$M��T7��0r4�|>����Ǽ��x/h0g@�~ǃH���T�]�������;�L�gc��,ty�λ���D�e��&��d}!l��48�M&���!:>m�D=Y�!yNyG��B�8�b�i���R�roj>� �-x����B��c!��[(3���~]�p�̄7���ĄЅ	ט����H�8%�X���%��cYjT�A>��p����@PW�W��B�������*���~/~Y>�o��b������~�{���|�M��b�1�b�ϸ/�d�'�^l~\�l�Y��=�����g���G?��3n�}<���~3>���/����x���c��^�߷]����"���m�e����-���v��_��/���㺏q�6��݌������[�)_l��������8�_��X{�jx�����Q��o����w���D}/�d7�e7�ԋM�vS����~g�2�ʦ�F=�%(�{|�iP���|���73䏍�^�fxƸ۵�h�:�e�cr�Ã;�_���{L�b\+F����~����c�[�������[b9}����K�Jj��?�t�JeǷPO��R�BQ���7�⃱�z��%���������6����u�?؏�%m�����5���Ώ�7��.�����|^��F��aһ��8-�[b}4'mӼ�~�[�a�z��G��yn�ۼ!n�6bƏ��v�?ޥ_7�G[��U��b���6מu��?��z8�W�Ub:�n������1��`��{��?����?�����_��ʛz��>�*��$^p�0�l�R:]p^�~2�?O�e>�`���{�J�9�,�@���4���%�|�͘�e>����t�^!�u��	P���h[��Y�+�̾nh��K|�(�g�]�}�\���=��`ץ�4���??�֏�p~?�y�o���r�4��iu��O�ŷ=X<?�=���g�ݼ�Ϩ���o�'^/��cn.6�\����n�߷A�s3n�巋���f���`˷)����>������}�C��M#���Ώ	4j;��^Y��Ϗ�56���Dsq���i�<�89�?&*���_S{m�R������?z�&��M�P���\~�pk&��iԱ�{o�\Ū�>��P�)�B����|*��+�Z�dp}� ��Z�c~��p.g�9?>s_����J�����;���o���@M��ˁ�&��;���n?{��p��7��p�?�5��q�uG޺����ȕ~��g^���W/�.�/�����!�x�"���/���E��u�h���8_drS�.�ojxיA�$�{l}����H�p�7 ���x�v��~y���;����ߺ�������۰�\�����߾��纴/2�+.ǋ������e�{3�\ʥ?3e`��ֆ�<�?����i�ȍ���'���ysH_doG��3o��2ܒ���"���F�����g��"�ߊ�u��sS�__z�w��o}V�?���!�oG��n�@9���E|D�{��`D���ɽ�C�{g�UW��ޏ������Ϳtw��fW\�t<�c~c����Ϟ���^�_{���7���n6֝�x�x�{�E�@�&��.��󋄿��bǥ�~���Ӌ, n%bx;�|L�m�a�!��al_�b��q�w/�_>�>Yq/�}Xe�-�C�"�	ټ}�eb_��-yO^����8amr����ancni3|��@�W�LQ	k|���2��!�G�'��E܇<����V=�G˙�y���|�{gᷖ��
4d�=<�G�	��Ox4d{��YP8�h��p����T�X�����݊C�����S�ڃL���F��ƴ�����yyXsc�Ok� *I8�8=�I�Ͷ��QA�JQZr��FC7����:��h�9+� @���Z��.�u�0|;�O[�т���Ĳ ��:��k;̴�����@UAԴI�SɖH�i��|�*����-�5��(cbO��f�<Ϥ o�6�@ =4�-�/"t[�bU�)^��x�=D�lA�S �} �M���M���8G��t�3Z�W(��<J�M���oA00�V�I%�<�Λ����g��B\���`�F�j��^����^��?��a�008B�����O-4��V[Ȝ�)��ܨ�%`�6� ��]u����*�������Ҩ�%�S�Ybyxz�PJ�&ܠh��զ����6����n������O�&;0�6nJ��� �}�,0\�}����K�Ë�F�@"� �WЈ@ �[֎@:eda���ۂ ��_���<ܺ|@<�R�> �^��Haȑ8� �D�N_�i�Ǥ���D�}#%��O�������-��Q>;�8��y_-A�V�ϴL��F*�+_����1�	��d.��m@N(���0�+��!$
�U	i�s?��Ёʴ ��O����V��ퟬ�y��%Tr��?�-f��$��Mth�R.�]Em} tR����%p����bg@�ުx @H=�bL���!|cC&P�� (�B�� �᭪�UK/�c��Ҫ��/�g
���B��ws�E����;�Z{�� ��rYZ_P�]An��f��P��Kf��������H��KS�<�'n�s*��
r���c5��|} %Y� � ?B�$��[�N�uA�P
���^f�ذ9��6@hSe�~�CuuA����>�y�)��'���~ �}_A��[$�,'R�}�"@#�7A0��0yoO�@�	�NA���N���,"`j'�d�٫y�l_�&�<S��;}��I�B�q'l_ ���rup�o��WA^�n�e'� ��F�W�zC�0�6$�F�u�8��dx�z�8�o��
��@�����=�*��ď���~"�_�ߋJ@����C�_�"mB%��.s;�b��{�B� �W>�������'�*��e/�$�W+�_<�k�g`*��Qx�-��Lߨ�D> ɭ�,��Ap1#�ِ�+p1N�a�x@ 4�� w1�[�̍��Uy?�eb�`��Y;lOe�|�.��ƃ��p3g䤹�<�u��xlB� /)Uo�6��÷ ����h���t+_Ah	�[�B�o�
B��/�)د�A�SyB^{m�|�t(ǕK�9�;nG� �/�Oa�v�&%��ڃMjtluG)TA�l�!A�*VwAN�#]�I���o���� �C��A�,ȏ�� �Ԡ���|���#r�>���9��nN&̀� �:�0|.�� �����	�X��i���fA���4VMݩ�Q8��-���u�Χ��/U<5�c��>q�$4!���5��'�����Y;p�i$A��w,��b{� o|�w/���Ɔ�����-A���Ԯ�9�8L�A��v��Z�1���]� |�}� S��`���" ���a"o��k�&��Z�A�;�����;꭪!�!^6����C��(o1��6pQ2J#١��Z�y!,2�^�Ďud�`J��	�jE�A~�1x�'M�uNa�$��KI
���Z�F%��F����� L�āK�Rx%����+L���Q��Al���|B��G���:�ċ�2'�^����vH�>�aѕ�Wh>Pi-���W��@�{>p&�7'U�^��S�{|Z �	�UC	����o�V�YY��域4������#ȭo�2r �gZA(�¬X5@���K8߈�l�f�T��g���]����AD������ ���J��r��N w�����4� o��eAhՎ���q�&�M��Q��<���I���P<(�v�� �	b%�c��jAx
�ډ�^8��ۭ9@:��I}�98k����s{�v^f����p���_ѷ�,h���9�=]��/j��0qW>'X���7a<�p�n~��^.mEA������ܜ��x�C7r�Oa9Y��j��	���$���D.ډ51;�¢�p#%�7��t�sᶹ6�(�|�\1�����vCߤ.u�7���~ämP��D�8q��
�j��\|����O�����WLtZL�W@#{��[��~�#���~a �D�"�>�PāQ`�� ��D(�f;��D�P]��7&mt"�c&����Ic��;-� �O��AH����8`�/��UR/�|�4"�����O�`1�����q��U�J�e�AP� ��#���-\���U���䫸� �ﻨU��֬ZO��$p=P�.yTs{=�_�K��!$1`R�/M��9Aޏ�!�m5�=
�-��=�jP9�ҢJX��u0Ư
�sa����iu�����W�#x\����q6�:♖��wZ? # #g��-^?��lA�\��3_�5�A��Q��G)k�jY�^��W k ���>��G�^�:x
�Nk�U'm�lh�����|DO�U�^Įi��\^3�B��\_��	5�5q�&Σ��Q�p(w'k��[g
k!�D���u�B4�^�Z4V'���ǧ��k�x�Ȃ�Z���I*�g1Pu���Z�{��3/k#ؾ6:ު����� L����X���bQmX��7����Mf��X�7�~�s_L�[��Z�U\�U\G�k#� �D<�M^A��̛�+���F�U�"�R�9	em�B�a��)��>��P6L�l~����V�B̼ L�D<�L����&�l�)�J�)�ӕ؞�&�Ȉ[��Z������)�;-LG�c��A����}8n^�\�*��@xz�[�J������A$� 9A���
BU�+��0�
��r򬭬��{�t�w	�8���t��[��`-h;��zA~�'����3�MAlA�Eܰ�c�MFAx��xȝ�� �)��nH��u�&�X��/.����Z`�4�(�Q��Y^��])>&:t�
��y#��c	(*]<�H��a�7����h�s�;n*l�J��,7x�7?�~���T�0��r�����͛�=���e��N���F�"-�=�<쉵C�;"����~BT���F��!�d" w�k�M��lO�BoOd��%sσ9�}���,N��� �k�	�W�����^�G.�����i��|�2^Q�������ĵaR�W[�|W��|�����7rO�Ǝb3[lo�jk�AU{#t30Q�-���q�X��A�J������}��P �V�c 	s�,��_�owL��.`�GAh�@�� 4tltZ js�17ӹa���O��U?̠�� A��߉Ȯ"�AYN�6��C��ԧn7Q<�7�ha�P�J�=nnw"�'X�6yDa}<HX�9�:8��r�;�B��%�>8���~p�%s�I�b��+_�H ?�^?Ń�6 �C-@>&��J<8^�/FI����m;}�(ţk��:�j���E����`'�jz<�D�h��
�r�2$���F�ώ���,y4$~��D��k���(��{4���g��=+����p�<A�b��A8�=�o��2�������<:rk�r��"Ҋ�^ǯaD��g|A�RA��t��zUG�X`_�9v7�Hռq"o����H���K�G�=F%��9��Ǩ*���!���;&"f�t �ņ�8��q�1qS)9��t��^�1'ZbN?؈
�ħ@D3~@��T����PU��E!���`�.�� �i,0�rg+R5a�Y��b�+�c!B�B|t�z3H}Z�7�B� ���Op�[4a�{WwT>&66��뵱u��_�^D � �C��Zr0|y�2��0rvn�'�T�B�Q��8B&��ۂ�8�i��Q��ѕ�_����%� zĐ�F���*�I�k "���tG�n��C�P�{�=�˂uA�=��hRA�MWF��S}6	�%ApN�Lj@~#���� <�D�f0~5�z�+A��y���i~#-q�#g�q;���q�����Q� ?��V=�a�5.7 _k��/�	��$)� ������W�-���Ed��H�:�BU��P?��qC������"����d�iA�Cy���/��UA�f
r��giI�A>k����|�CE��\��r6�%���_�\m�"�˲�>j[�1�ƃ_� �Nn���Y9��AR6I-A��>fvl���
�_��Z,}+�A��OA>�s44�@P� 7�%t�U%EL�"F� ��� ~69ǧe�7?���Bb�Y1U,��� �rGDq��Y_��$�MA|
����k��rv��$6e�`sx}�}���uOȻc"U�vru�Zu6t��� ����'ظ��9Ao�d�I�ħ`:(�"n����gZ90�&B*
B�pϗ<7�	���P����yUG΢�\8��Ŷ\�S+r��_����=`�/�	�*�p�]���dxA(�����-���yt2�4�[*��d�@	%zY���i�v[���aWn0���B�'�p��K;7>EGd�z@��N��N��)�[nd	�o����G�IM���KF���/LF�򰑂��t�c�I� ֞�*h1c���KƦ�`'�� :����c"�@&��#�2���^Ddj	�xY�H�L\%�_��e��'�	>�$�� �0	fhA0|Z�|*hY��`�M�Fe"�5��6A!{��FAX��8�����(���xŃ��>8 �3�A��gb�t�RI�ensp!&���Q���۬]-�
.��E��F��A^���0�CW��u� ��Y�*�ϮDT1�����PF�;�����σ;��w�5�}a��e��μ _;*	�kߐP �W�ӂU�:�aP�)�*��"#�g��8�!��xQ���fA>�:r����tD>�m�!�q�L�xв�����8�?�w%c탩�"�t��i��o�����#���P�P`�0��0�� ��xy�(X�ܻ��_��X�3��~�!�ݻC�C嗂|��v<A�3ʼF;U����D `A�8B<�|i��΄A��Vz^�ٶF����C��3� �t��w/-���'��d/1������	<�@b��a���)��	�p-Ƚ���AXm�|� �
��|�)]���p����D��܇�=^�	� ��pA��i��|�.��7?�>��Џ'��`�����t�(
���d�"P���3>A�=�&��6�OEC��f�� ��k�ϙa>2����A�*�8����a� 4N��U� M� �a� v44�
B���
�ѢgB�$����A0V��P�$P�C{k@ ><�=d�>�XkAX	֕�� �(=� [�,�p�.�v�^��}�E:89�o��S2����?�6�@>��F�[Bu����9��	iS�ŋ]�������`�����}�`y���bw�`�����/�wo��;|�zh���/v#�>؏����l�{o�[xNx�]���ݳ�6���zw�]�M��b�_g[���W8�%��'][?�wof.v��>XG��x���~�ͺ�c�������۷�w��`��/_�����:��̷>X�>ئ}p���7��:�mv��J*]lqn��_,~|����`����]���}��wo�����sa?���ϱ�C���1>�e<�G�a�������7O���x����%�jtΙ�9W����k�'�������~���������}8�/6h_>1_u�WN�b7��b?�e|��a;��}��:��o\y�/����u<?X�o|�;>X��Vc�|���ƺ���%��������S���`���Q_��}3�^p�{cu���!<�љ�?4n��}�ݴ�O��������2����	+����\����z~�a��3o�ϭ縱̻���ЍN��~�Ϸ?�Lmq׏ׯr�'��5~{�$j��K�w�<w"z��χ��3����?≟A{I�C������ 7����!�׵̰��=�?ڳ�D�����{�����P}&�������M|��؛}�I��u5���#̣�_��,!��!��(���+=���+��u���9����e.�O��/z�L���i���ό��v�s��1A7X�c o���gѻ������?����x��?�5���{^��k�?�Fb��|����ҟ8V� ~{���.M��.U�q�c����"͐�Ə����!�|�E���e0�C�@�����E������M1�C�����{��"�i�r�'/�n�_��o�l�����9�G�����ކ����!�{G��}n��3�!W,�EP�J���'���Mr~��/M|�],���i�">V��|���T����^�H�[��L7�����c���q������b��Zu�[���⾈ϔq��||�~� ^�gӸ�����x��]^d- ��%��C�ϦO��������S/2�d̝�}dN�׼�1Ht/9��� �����ƺ�2/�cl5��ս/֕�~���t��k�L)~yC����F�"���5n��5\�;�f�H����h���gm|�F9��}]�	G���u�U�3�O��}V��#�h2n������}��{��ݗ�Yn�����`��ὼc��G�-|i������{X<c�\��i6S�4_=�y��$X}b���׸��L	�T�?d�Ȍ�#<��׋�@}Іq���P9Ά`��(4���g���t���-[n�H��"e���.��F�{)yP��~o�-�����'r�E|�<Ϳ�t�3|$��lG|�G�O��9�|����c�#��"{��\7�x
l��.	���Iy��:7���"���E,A~�ߞ�M�<�M�z���_oQ͡����֐���yT� �j��u���j�k2�A��]1�GPAA���h*AhUJ�
�qAD���
�����ZAK����1�T`ܵ �:�t$O�w|c��X�ȩ��� �����Hu���8a:�PZ-ĪB٬�	���DG"���b
�Al*�cb��/"�x'������c�y,Xݘ��@�[��=�@�{#Ş �	���:7��JZA|����"�#qB� �� �"�����x��DwA��D��&V�	*��'ĕ9�y � �ǉ��J�AY��)40�'���c�\�����8�:�D����&�y�a�`�m30L&8�ՋX&2r���NL0a7�����փ�^t�y\� ��l�����,s�\��00�y��������~\H�n��<\S���N+%@ ��(�t6ȧau�H��սK��� �ml�X������7�FLr�H
��`��[���N�s;8���dF�1^+�V���!A(~���n��|�h��a�������ၾ��� .,� �0tkə��	>*AXʩ��i5�_ŋ ��V�,�����/7V�Yj��Z+�����L�/
bKp#uh���� �MvM��y%m�"CA�D�/rM;tj�']����Y�~
H�h��n�v�2?Ak��A; /Ȇ\g�v�>���3A�F������]��U�r��$��E4^c� 7C�|ޟ�-xq��)߁����>��/���N�%@��A���ݳ��q�b�Mؐ�U��(k� Vbz�Z'1@����]5(�U�S:��u��	r�*c�CET���:!�1�^T&�r�PfTM��
¬�Ц(�Gaל |�� �ou�@ޮ _Ԃh�*Ah	A|
�=���EZ��Jr@�ٵTQ�$A�L���@ �]K��>����͝.�܏.�D�ŉMl�4z'�� ߨW_�I���DȂ���|� {�("�������_�0a&����R� ��Bbm�7�-Z������@�-���YUZ��z�5�:~�$�=kA��~0�7������oPw��Mi�� o��{���ۭ�A"&vu��\#�ݾ��� ��Z��b�T�o<��/�#�DǺM*�^
?�`�KI̐�t�>�^�%��Hܻؾ�+/�E����(��{��F�D��G�$z�ڨ3{\��u
�wj����o��y�)��8=ُ9ф��nA�����~H^\~$V�����=���	��N�x9i�����N�y��S�P�����ӻ~��$&*K���K;����'�cR%���v��5�@Ū����}�X��	�o���5�d��,����E��2c�V�6>�o~���A�V*���ڕ��܂�Ut|ұ^KSe��E��6� ��Oy6؜��A��Gw4p,�\~��EL��+A��B��V��D��C��A���zQJ^�L_�a�u�p
�v�x
2S�ܡ��J[�S�Z䛟��\Q����/����;|A0
2����zȫ���)�U��W��yA���C�H��V����XA0����������^-�o��H�oħ0&F��#�MLA�TՂP��5m�r|L0V��Wu� � S�1��#]K��1A9.��0p�s�M�����A���wWy�4���N0Wʋ���X��p��٫�YSs{�I��EweuL���ʱ0Y� �n~4�1 .p��Y�-L_�`�|s-�k��a`����'+1�CDicCT��A�zሺ��7�N�
T@���l::>9�BN�d�}�4b�x�2a��I�ذ䂼�AU#ت�1�G����%��D��y�0�~a��P�v��Pyɤ9%�Q"\q*$.]�q�3��#7�n��rc$�Gq�;�x�qh����!�l�Cg�@(@|���|<������,m�,!<�;CA�Mra}�� ���7i��|�q-��|�)-��Rz����z>p�B���FT���0
�����w'�u���� ?㓏�^�lý�P���n�P��޶ >�_�[���QʂN���wv�dr�3;��١�TJZ(�A%J���V�D�������!!c��;�bK@�m�^gc�v�<κk ��dv�����������?K� �ѥ�`� �k��er>({�@z� wj� `0�98&�����+��a:>����wN��	�-��_���S`�����i��%� Ah�	�dA�*NF��]fm~�&m"kNY����u��|�3qt>t�'y��L� ����W��s�h@�{�s! W�����]����h��q_+�/�&/��٘��%s#�G,��p}v���ܜ
�C遲�S�ު���ƭ� ~6ԏa��P6�J���(}���F$j	�g#�qjی���_<X��q�\j�A�P��A�c�BU�1iS2_�m��P{��	�A�8�:���\eMF���0_���HE�)�88�ٓ1�z�>��I�q���H��	�LKd��yp��c�D��3�C᱂�<6�A�o��z{��3A���������~���r+�\���0�aDA|�[u=8�[N��g�O���z�= �� �:����X��UT�;�끌٢T��-# �C����k�z7$�7׫�vK/ T�!\������B���(A�}C@� �=�WC
C%o�7�o���j�v]y����G����A�=]�����	�t�.�6��o��{w���p��.��An1��*�[�#���cQ<������S���y�uvGE�8��7A��	��0Ȍ��L`���[5�/�r�}�(EmLܕr� ��k���Z�o��K[������kjm�0)��(K����^�0|��/eA�jq�&Ts�k'��+�І5�&O��� ������ŋ�r�~��р ��y`:N;����x�/�①���&�k-?�^� �"]��&��c!�c1�~m\��z�jQ��mk#�Z��9��!FY����	h8/�E�� ч���D1H+pٸw�Ŋ��P���H�Z�0�L���ΎDT� �6��Ɇ?;�\"E��)�Dt� L�I)����p%��l(.���ơ�98�(�_<�����A�oA؊����݅�LB�0a��t/MG@�1E-^mi:��[ܕ��X2�� �ݝ��0�� }d?��\���u��B
��p3l&2om� ���)��R!���n���s[�GLME8�)�}�º�C\��ӡ�An1�,��	�%`7�����N���Mv����n�mmݼ;�O��z%:&�_E�vdA�C}�5�����M�oA�=n�aZu���ow�F�J��� 7|�c�"�7����B��~|� �6��[��k4���~,S��!� ?
3����$^˨2ً��XhBʆ�Ө�P/\�iW����Љ!7p��'��
���Ȉ+?�+1����е!�Z9<"H��>��o\��#�c��(k5�:�� �����O]�����XH����7��dB�0��{�,go�4o^Imt�\2�}`Mxg(3m��
�(ܸ1�;a17|ߢ9�/���;\�����@ � tmt��L�>ʻ68�'͂0���X/���Ng�D��Aw}L�x	�� ���9��dA(^�����'�4a�r¤i����C��>@bw"S!�GQ~���@y]|�C3t�6%�Vӑ�cLh� ܇��AH����f;jO��L�����n�qi��{wA���.�AP� ��'ل���c�(�3@���{�}Uޞ
�a<�r�����]����Z!�QV��ZA�)ă��` � ��|;/�V�X�?(}}�s��$�^H��5�_lp���h�޻h�� �{��Eh��M�p�>� �0Řɧ����ҧh0�� |����;&_I��	D+�!�!>��zt�䣰��wX�׏,�#�S�W/� L���g
ARyA�&m�X�΂���І����0��,�ʕ�7�NK�A�%�ݨ�X��0�=3��Oֻv�B� �Ɓ}G��6p�S��UA�*n2��Ȃ`����qQ0�;���L@Y w�g�9p Zd�����Ъ�s���U�F�+��� y{m�V��=YH��d��`���L?��:�k�D�	���� ��b=XtV��Ą�X�U��CA��V�� ����S���C�suV�u`�׏&�2���ѷ����S� �yA^��PA���=1L6v���8B,��k�/6�oc�bI^�08V�c5@g$Kf�ĈD�lU;w�w�X	��Ep���aU�+�2����Zڅ�ہ�H���kDA�Ǥ���\c�͏RT-?g�� 2|G"$� LIo;^ZriJ�N��� W��cRA~ZY�qX{R\�k�����^��#z�K�FN>8�g
5��!X�|��3�	󁂏 �V�|;��n��n��.� ���YA��(UE&UQ�y%�+�}���&l��|�%)���I��l�X(ȿ�!�R�������E� ���	�c�l �̎�͂���A>���E���l�$�.-J<5��&�+=�/=�a�R;|L� ?K+����A/�U���A�(�O��M��Q����}� �ӂ ��N����/�� ��O!T+�(U���fh U@�{
Z���ޞPOJr=���	��SE��E*ȿqN����m�|��N���Ή�uA�="��$ւ0�&��ypIN�.b�}Q.�'n�@ϓ	�`'x��T��[݂���AB�0k�m^-'�|s���MY��PsmD�'�s#@+��[�ܸ�,��&�`UˍD��~�����M�C��
��S�E��ߐ�ˍ����u�9�CP��l� �g��3���p��X6��P�{dA����ܰ�z!/34%KM~N�#����`���R�.�E��gBi"�� �19r��+��`|͚���ZC�� 	�^A0C�x�<��A�bU8��Q��P�%%/��@ĭ�����A�c��|���$j�7e�<`�;8	�3M������D��y��	A��}�	r#*��A>��2�A�!�֡ Uq�����y@�W��!�y���f��@�l�BAn��=��5�|m�_�a�(����C�:L���i�Ӥ��'�'LA�ATH�F�4�ZA~�T����|J�ʂ\�i`z��4��
���/ߺ����iǏ��;�>/v}/�t�bw�[�Q����C%����y8�^�!�yC�� �d8��t:vM�c?tJ1,fO?�>K�����ڡ�#g����L�0,\&�@������U�܍�u�� �� �"��c-����A�&dK�2MP�	BU'H���L��z����^��6#���B�>�;��q���!��ħ`�'�ZAŠ�c��8E�bŋ�8I��`}��
��+#�!��B�MAn����%� 4�B�� t��>�,�"Uj����6n�M3�!�{6��
���=J�g#�Hl����(cU�7!��+|�_$S�	��=�ct,�������o�Y	�v�X2�����k;�FAn�����@^<���C�r	�˓H�=d��6�����)e!�� ���%
�z�Z�����a�ZV䃤B�N�4�?� �Ʌ��z�	��:H�Ǆ~<`�-e���HAlB\,����P<�~�C�ä��{FBA���z��	i�ܰ�]E����Z���ύכ�`���\��z����b�͗�`�i�`��{��>�a�oJ��Ώ���/�~[{�n����5�[���vô>؏��!��,﮺l�ݛ���m�&�P�?�r��/?���4l�Mc�.�1�.���n���h�~y�?ۯ��Ӌ݌����R|0~G�[�2H\l�������v���C�u��?��:߫�+�9`w��`u��o\����1>�~,�����c���;n&�ł�j�{��X�`��·vm>�/��|�˛��d6�������^}��>XG���e�6��x^F����7���n>�����x�b�G���zX�'���q-��{_��^~0έ�iK�����A[�.����_������+��U6����`ܨ�|r&�>��C��T������LJ�J�zv�'/��}���_�\΀�������V>nr����=�����������'K�`1��=�J�hD�s@�i�{l�i��-��5y��_͵O{n�zQ(�����P�m]i�[�s3�7�Rg�|8��O��"��u�?>����瑼�����}�����I��̸+��i�������?��ϓ���T�T���K�R��g��y3���|f�i��Ѡa)ǝݱM��z{����|7�/��I��;���0�
��n��l^��������n$�������~%^��?�}�5y�p�f�!�+���{/�z�H�����>�C�s#�!������Y��ڎ��uGǋG�Q��Ƚ*x��\�E�K�k/�[7��Eҿ�2 ���ߺ����ߐ��X9�昼�h@�VZ���>0��������Ǒ�6�\�:������ ��l���8�H:rc�.b�5��o���?�3�z��4/���">z�ݽ��[�ٽ������C��׼$s/��܄�lG|�
�3>�?�;���C���L�3����w�g?���u���Ч7G�>�2 ��ł�Z�#{�����!��sQ�>w�q�������ZW4���}8��R'�!������4��LoՏ/s<��yO�	�Jz�!�ܸ���s���>Zv��{��=�">2���	��h>�G�}Wt��}����=&��>@��x����E�/"}�
��J�.dZ��{w����W6_/��ɨ�C��omo��>�e�/�f��C,۹{��y��E�$2�J|�.2�8���`$��'���7au;��}l�i�C�����<���kQ	}j��)0��� ��.�Z��F�\A~i'�U��I�7�,�{��L<A��6�;�"��&l`�h�:mu�ׄ�<GE�%���Z�}Q{�-	�h�Rq������_C��m�<.�u𗴎<����:�g�n咢�(8�:��y��:��|%�냩C�E�C�a��6����2hc�`��m$�i)V�<H��
�P4ʀV�/^Dn��G�	��Vjڀ0kxX��k�H�G�i���M��֤�a�0@Ah���3�=����[�*���A���b˴@�[������퟽�Ua���y��P���d!V����hA<R��(LT�����B���^	�`s6��eU=��m�Fױ�J�`�lyTBug�m�I�ۣ2��"R�������C`Xn�����X�� P��,d���ז��i�h�l�����F!��*��!p�4u6ʂ�rc�W;���q~�X�0��
cu(е'P���v@l�DU�
���C ��P��nv�YtjW��~	�<"� �葁�aF�С _mBh�p�S��mAnW����������7,���2uR��e��K���a"-� �.��U��[���tt�
r�7d�
���dAn�d�=>�wdvr�ħ<W��&�0|������C9c�0�;4H:%{'D]���>An��-,"<�ĺ �ޖ��Ѐ`x�0\��Y�e���?�f� �R�^��ઃ<!�S=P����	A0C9��	<�+b�M�	=�boE��f�s�^�ύϞX��L̉�N�#gw�j������$[�"6��[{���o~a`.���<A���� ��k!c�B"��������$�m_��e9|�����8�CH���r}C�� T;C�*�z}�� "A�����N���q�׋xߠ�*X��	�5	��zńKlh}�c@��ԛ{`#U"D^�||cЩ��dK=9����C��0QFfG�M�L-����	Ap��|� �N��r��A.� O[��7E5����`�)��Na;�:SM�ɚ/�;g�QQ`/@n}�Ӽ^���t$ �_���䚸#R~^� _E�,4�x@�14R��.�ȷH���œBa4������"���E��*ܝ��A)ȷ��|cP��x9v�#�S���_�>H	0:��A�[���8���|�0�d�c?Al/0e�1L��%��8�+�N� _a�X�L��A>`���"=�r����/Nhj�Vr��Z;&�g��� wj��Ĉ��� X����B%�t��
#ȗ9A�Vۚ��ˬ����
����C>9!n�8���>x2/s{��Z��_��5��H.�Egc[��ִ�����6&���N���N� w�����&mO?%S_c�o��	BC��&��#�^A^���� �R�q<m#��@Goՠ[ ��+���ceA��2�d*�+��w�Ъ	�$�8X��ڑ�w:#L�	t$�	9�=e����� �ʒ�cu�I+A�g
�,�_���t���p�|#�@uNf���|�K#��0���|��&uq=n�y�ì,B��vTRj��Y�i��U�gbY`s�`�B~��A��5q/M�{�V��?yU��*Eҋo�j'ծK����Xf~R^�i��AS��_�0 :�rf����{ߞ
bY�@�w��%��ŏ��GA���s��r糶'���!A~0;��
�S��U<�w�\Q��3QA��M�����uH�o��F�A�+���%���е�-���� o{�g���g5'H���� ��	J�9A�T���k� t�#���[8��+�'*�p5?r����º-��G�'|?4)�T�|�=�I����r57|̹A�67����F]F��1� wBY8.����sn6Φq�����pA���.)B�� ��~��L����1r��^��@AX$��v㿘f(q�-S4~1'fZ�Ҹ o�\���L��h��*rn� �(�=�2&xꠇ���{��T��S�x.�rb�h�E�������w�
�-x�⩄�:Ѐ��䗍�A � w;׃ۇU9لP<���mAޏ�|D�L�K~4^�ҴL�y����q��l/ȗr�_�Ɔ��(˻(&T���'����X���aL4D��~��{��p�(�w�A�P���?_y����P��׎��aB�� _�W�i��]� tZ�e� _��^au�B]�wG�8�Z�GrT����u\�����U'z!_��\��F�b����Z('��B������ٳ/�λv�*�k?A�&؇��m� �xXU��9DA~����a�/D��_ۏx�N�-��0k�"f�M����@���^tm(�V(��~�|bQ�F[�*�e��m�M�� ���/۫�ܳZ;]�d1�^݈�H��8zZ1�>�@��ݯ<r��	o/F�k�	{/G�?�D>J�l����2%�$��+��	YˢNF%h��BK����4د�ф����F]���^i
�E��U�7Ρ=�7��|S����I�M�I��*u,@p���䝦=�_�����AB� _����A��
b�[9YG��[�W�!So3}7�O�#�'�/@nW�� �Zn�vC��f����mF��-�������4t��ͦ_X\���r�������ٶ\w;��wAު��T�Ө=��?L6�X�T�	���= ߽|�=�m��7�Y+�7!�7��ľvSn@��ڿ�B�y�ł0����G���w���P��[�������!�ʅ`sv�T���Q<[M����Z	BU7n�`0ij{{Q*P�V�׿1@ᾣ�2g�|1�G_EB�p_�,��Q��~�Mq�p6������7�w 6Jj���p�ЪT�����|�xA��@�Nh1��P�3��&���X!��`�N��t:�� �cSn@[��ê�V�&ǃ�8A>V��m`�%d�ƃ�`^fA�!�	r_N��{��ܸǃ�!A>a�N'85A*�����ގw��|�%���4x���њ�An��QԲ�>|�ᒽ2ͽ�A�Qd��FGC�V���^�o�T �7ߞ
B�ɂ��A�����y�j��
rˤM ��Z+��"���� L���8�n���$�K��G|c��9����_�0k��]�>��cҘ��1��|��<��8%S;q����B̀����,-e�ʭ�S���!$�X�"������`}��b���Y�Ba�<�&V`D/�̖��7�:��c�μ��Dμ�K{7<�͵:FtCg8(�-����Q���LG �� o�@�� �
��VA~�&Xt,ҁhAp�98��~yj���ȱ|�]~q�H8��f �I� �ZrX	� 
�Jl�j'⍓�O� oUf6F�Mu��c�EPr� T����8r�'nqh�����``u0�Z��<T�*���P�K[>��
��8���;T�H�0 ��_��I�Ţ��a����)��N�*1�� ���A,����m��U�T,���-��V� �z_��!ļ��QN���ٶ���G&���	APfopaK��?��y侜 (�w���
~�U�׾c[#����O�츚Ɏ����w4���H� ��S��`�T�cZP��D��#�~��*G����>Br�+�|g(ȏ��ȟ���̉8_�av��� <�3'b��{�sa*L�K	b��3��H����Wb�q+�aB�
[ OH��	�YP���0&]1��N1a�1	�Q�F�2>Z���l�u�H/�[�;"ɌKA~V�£��y�Q�9�a��8@����cM�z�=rnZ��ҏEK��6vs��A�x��1�1�7eX�GbEׁ�pț�7M���
�������f2���Q��*/"I.�g? ���%h2n����;	Q��e����nAXN�-k��i� ?�ȃs߂����ɟ�S�p�z!x<6��`���U]+U=�_���<.:��Dσ3�� Md�C��P�~��/�O�о������)��V�|�+ȿ�=��^Ht9�iT�n�]AnN�OA(��-_���-?<����"��N�M�  m~Q�y�vЪ:���B��;U�����T�pSvx�R��EB��D����������D�#��b�����(Aj~<�P�O���		Bo���b�������g9c��-v��BY�w���. $��Ϟ�)��N���
�<�D$� �� ����'2]��5bŗ�q�&�WdX���3�~&��C)ȗ���X�/�����~qEfj� �,j���$5�Yȶ87���gw�Bu��6w`�0�6<�&�]gC��lĜ�����雐�F����� ��#��P	P�i�a��8��/{(��+��'_�?�Nȋ�=��;��1;�DD�V!���!�I�6����[ʓ�t9�H	��-!��U�I����/U=`�>��d9�=`�; T��� Vysu)�/���}��W����f9�f����ύs�X�b��C���	0����ޘ���>U�{z�{����8��I΋�K�s����^�ዡZ���t��X�v�I.6�<�
�ww�_���̵���ŏ�B��
���j^�ޮ~0��v�:>�F�����������w���X��>�b���߽�,���ӥ����1���|����ڸ;�Ʊ1�L��&�hܭ��Vgy�u�(�~�D���9=n��Œcc�f]�w6�����`�ؠݘ?���yt_��{�i_m5�m ��r��ݸ���z���:��߶���l�u�Z?�D�}���R���h\7���Ǐk}AM%>���ߕ��W��>��%�̛�x��w�_��L���{ex������wg=۸۟_??�~Ӎ���4]���q9?`�A43�Y4�x2����37��i��s��u����v����a��F�a�����O^����G���J7��~f6ֳ�'Q%���A6��p�}��؞�(��Ł*����}����uw�w��]��>����F}����z��cr�9���Jr(^	����f������e����g��5��ߍ�?����0�����e\+���y���.����������+�q]ZG\H�=.��n���\��CF�".U�ay|�n�����e��C6���l��%��������?��r\~��&��ǿ�߭��\�������ݢ�!˅��,G�O�r��~#�����}�����.u�/���>��%����#s8��OGs���qS�����c�FÅ��5�/����}: m?���q������;#PûU�C�������|6}�:����yv��s���Å��z��8�����Xn[��!�޿b���Vbn�V������������g�'=��]����|�~�x����Iྈ�y]���3�m�.�E|-X�g�B��Y��{p�؋,G��˿��:��u	���o��#;��$�"�����3�W�=���{���L��=}��{�s/y{�t�����x�J�j<>���Z�W��x��f��to��x���Wt��>�b��^�%a�C��a,﯀m�%o���C��"��Db����I�?yi�^d�#�6��>Ib}φr�u�ҽ}����7s����p��I��,��v˖�7�EP�$��8��$���<����|�?ݭ��Ɲ�����@N ������5�l	g�X�����[�>O?��/���u�3y|n]�4B�d*�4�B�:k^M�B��ٯ�*��oȗ?�䁽��@�)�OB��嬶�lg	���B�(����rxÍ� �3�5��B�V%�"�\[;~E-2��xW�����~�$��^�Ԝ��N눰hw��FWm���n[����xA�|}c�t
�w��V�$^L�+�N��}P� m#_� Ԟ�łX<x6�`?�x��`�6�_���.��hق���-����I�9ay�I��ᩀ�%'� ����ʂm�'X�D�B��;k��`s&�V�D�ocU����{�Qp�0�&2��D�g+bx�����b\�`hm�A?.$�
���J�_\�2n����Y�ڨ�;�/���~Z`<� T�-��UZ��H/P�7�Ե6�Vt�mP��ݱ�CԵ����|���`m��==ү ��M[�!��6�x�U� ��ɯ�0�6RZa�=Q�>�)�c {��֭}v����l�NA&fbApj�- �ӊ��!Z� ��<2���m^�JwL\-A�(�B[�';�F�ꖈЯP�"�*��Aؖ��/�-����n�Ъ�ᳩK-��j�v�!Ҵ��SP�i�˂��P��7������8P2�{�Qx�y[� rN�An:
Z��"������� ɡ���?`�YumO�Apӵ��9TZ�|
�]�w@�E0��Q�l�o<{Gso n��Qھa�
��N&A����Q�|���\�
��{��|����n:�^����UU����âq��/b�-�C�/���zz�����T�֞�MG��%��\A ʨ������n�-y������B =�b��`&� �"
�Bx�
�/B�O=	� XH�;|A~�Qw�^��1V���f�/�}��h+�z�D+���������*� /"s�o� ���C�}CL�ox
}���!\�`�,BH���A��#kӱ���7�����N���]�h� �j@^��L�~��r�����~�$���
��
h�Td	Z�3��h�'a�%���D/"C�'(�z�M�S���
�`�+O!ߺ'�y~��)x�=��[������NG��)�0�rD�P�EA�_d���QT䣷7�0��;x�R�� �������ƃs�Q�u_2����.7ƃ�A p2_P�N��l��a<��i����ŧ��&�m�xp2/ȷ5�A�i4\�R@�(<%�G��o��킼��D�y4p�
Bw4�a�B� �5t��D����������Ԏ��.st����xZ��<�<~������"���5��=�׀�����6g�|�� A�8qc�ٮ Ho�A~hY�������	M�,ӄk-���-� ?�s�X��� �"6,���-�s�	n��ċ�DY�/7)�a�X ~)�u��R: -��D9���jS��XA���>�X8�k��hm2��7$��&�`S$�|7c��XC	3moL���Ar;�7{��A�2�
=�cEl�F���G�L`>j��-�em������� �w��X n
p�y�F�@�jP<}��� W� V"�%���~�q�;J>��:�*���q �V�^�C���qpli��~� ���O� ����q&���k���G����gC���P� ċ� Z�S��A�h�����p>���W����p;��ۂ:�g��2��5;�GAn�&	�f� w1
�v*�rx.�N�d<�� ���g�w�� ώ�����Im�J�����l�E����QH?�m�Y�n�\970spZ���9@[S9����x�eMh�i��1�����a"O�K2^��}NU͉U� o�yܽ�y���N�������:�R5�6�~�;�1��1C���)����@�$�-�̹�*Cn?�Z���P���4���q6�#'��6ΐ���mN>�NF�̍�-A9G�0�6Ng��.�
��� ؜��� ��Ѥ�� ̴ Se�d��	g^�;H3�1���O��)�g'�Dg��j�����m� ?��`_��W�F�+q8aH5a�P��b����d3��eCa������)��?��a�{{�<^��D�Z�˅]!���C F[� �+�^�Vh�?��}-0���3����
	�E��"^�Sr�wM��ʂ r���CݷH��<\��/W3xj@C�q��l[˄/��h@��4���j��\G)u{�&���j��_���-��a5Z�i���w�P��AL+��#i1scux�Z�݅]:FZ��C�� ݈���v�``D��:�w��k`�)�5�#)�w �t����__�� ��ɩŬ�G��}����r��O0/�h��+��5��	��"�� X�r~��'��
k"Tm1�-��ȵ�Υ���B�]A������,�H����Ea�T%M�qC�6g�`C��1����%`�~H�o�c���o��_�B�q�q�$�w�K\�r�+�(r.�������CA>Lbb��e�`'ѷ+6�⾣ �=�x� X����J���:��u]5�����4./B�� >�J�<&Vb�,�M���*V��ه�,�$��b� �t��C�s�����(�}�� ��`�������(,����Bd���)/"���2Q/�'	�I����پ�'���S~״H�
�S���>�n����]�ᠱ �=c�w�)��k��{�u����n`�V3�ºܻ��_�� m��;����f̼ _X�w@Y����)�O�>m3uz3$S�c(����r`���8�U� gR��� 7�{�n� o���w(|&ȷ�E���� ������N\��	��X��"4�~hO�<��֦���. /Bg� o/����k��oh�l����J&�Br� ?���)e�;��q�!������8
�8o��ب�И��ZA��jV�"��a�n�)#-~11�6����)��^����
�ҕ���h�v���kc`��HnJ����A��)���y���W����B�3�E�;?��-�מ��|��3�rV+ACe�K�����fh� ���1q:��t���a� 8H������:zA(���P/�¬��^j�@(�0�2pa�=���ÿ?���M�D>ǛPFȭoЙ:��,$�T���磼	?A��I<˧U������OA�nr�.*�O��� w��9���a���Ne�����Y�a�
��ō�������/�CL)X�pX�E�o�@���J�;���qp�������-f��>� ��r�C�(ƽvn��t'0H8%�MG���Emj��T��T4?��9���BP{Ax
l\�|�+�|��X�ƁDA�"r��Q!ƀ��A��T�H2�\G��ɹ͋��EIp�$�O�bbKY
h^���3��W�)x	Q1��Wj��AA0CtYu�̧0&HV�U5����{A�����G]o��&[� ��~,�!� X�:�0ԑ����^A^�^��4
̓�O������*6������>O-����8$��8wAX�x��KS�C^�>M;$؜�c_��9A0�2����}� ?z��*p�%�0p`,��j#�>]���ڠq0��&�O�T��0��B�H?T�Ml$�yx� T"~1�"'rk�9M��'�|�V	�(��s��%A*�J�A%��	��`�� �Q�X��т0��A�ۭ�8&Z�mD�?S��]��!� ��s��2D���H>�b��� �Tc�-S>���^Gŗ�)d"�Z�.� ��)�Rj��]@��Y�fC<yA��
�|��ͲW��`P��&٦[�l`r�C�ou� �LA�c����P��|ٰa�'�IF�| ��C-�������9���G� U-ȗ9_̴�^GAx!;����貒Y3I��ݽmAn��Yěp�)���<�A~̐d�-��1� ��pA�'3pj�����k9��<�!g�3���"�Dƒ ?���ρ�1�ב^ZN���\���ۙ��ɉ�ǜ�,��`�.ܻ����d�����M���sI�!xKP�>������v�zmШ��Ϥ��8@�=0�7�r〽�#���"�E��ץ��Gf�ks��D��gp\~�\^���H����9��UV���2�x���� ߱f��$�_�Hl)3�Y��#�Q"�<�,/c"q�/�J�`P^:�v�P�o�ʽ�/��<~�r4!X�xy�T�Є�x{��	� 8����a�9H��5�IVуKЊ��!~"nka�ܕ���L<��yJh���y�m�y��A � ?��K�y�L�̓���x ��>d��VN�ם��E�/�F�O�CiA��D5�|
b���  �X{�P��r�x\�rӡݼ�b����T��|cp�hAh�N8A~4 �W��K=A���S� �|	8�,V#!��N�Q8-1&2gO��>�~�o��#�A>��̟�#���"NjN��p>��/�$���Ym+�ӿq<0V~���y � ���L�ȇ2/����"j��)A�q��<�yg��O�h�������@�3q�+�ų�A	g"Q� >�!7A�/y"j�,�0���͂�"�a0-p��q_�?�����P�� 1�Y8����Q�gC��l����:����k�/A,Q�0rx�u*�*�[�CᏳ�;9��؊�'�$w(O �EL�9���W5p�,ȝSA����4 Y؉�)��I�c��00�$�OBVB�\B�P��hׄل�	�}��<X��
'A<]��or��u��zhR	�#��EA~�v$v
��:�
.�Fo������ |B����>~�$�5���B�=��⃽a/�m������w�{Xz�K?|��_��� ��>�nl�6��Əw'��ݫ���}(>��o�,���_؏������߽����M$��ݹ|�����/6~b�� �Y���{��k_lqL~X>��sW�����m����7v3?^l<C�a_5�����;��߸qK���cL�ɏ`��n�����XW��b�6� ~�A��~0ڜq��^l>�"�Y�98���?���os�]�f_����y/�?؏�~��yG.vh?x,Q�z���Y~�������^�����k����������Zם�/X�� �'����$X{n�P��_p�;��z�����۽�O�Kgx�h��_��2��_�h�~���l��O��=��~�}�?���Ӟ����I���^>\�\���{��i��s}_��J�^���?���>�]�}���Ck|_���E=6GH�����^'~��f�}�u�?}�V~���3�����]�>]���s5L?�t#Ho�|�g��N�wl���I��;(����p�?��a�n�����?�t�����o�����+㪠��_��#����1�6㋼��t����T��=��Cn�ߋ���Eޝ��Q��3�!���� y�������o��!���E��s�C��{�)�Cn�׋��g����/���E�ߺ<�/�Z�?dy�����{����r�"��=�#���ؼ�/�_:���I��e�}���o��ާ��?���|W���z��n����!�"˾T�ˑ�3n]��?�f�!��~|�歱��^��f_�K����L�H8�}�n؍}�`_�{g���W2zy�k�H��F?��1��c����V"n��Eeu��މ|��=�����:4q�m�o���'紾�彜���E�w2|�g�����CLt�3�FޭЋ��L̝sձ_��:?�aG|u8�g��>2��pn�̋����@���^C���x˟��_������d��^����Zg�cթCw$浯�/"©=���A��	�c3V�1�A��߷D����  ��~y[~&���h`v�'�.� �����Ӧ���/(gJ��O�)����A�.�ﲛ6M���sAd����� �>@,m_�a��i$0m�6ȯ�� �\ �i�)Q���FQ`�C�tk$�(@ :�o��7+�-�!A^�ɖ�H�o���d��Cy�M�����
�i���R2���A~,Stmz���p�
L땘i2&(�9�A�m#�Q�W[\��b%rIF��C�C��-��@Z@�*��~	.��a��ks�_0|��^A+тc"6Z��^�=�w�*�?9�����A���\EҮ-�W��^�D oK$䝖�iԽm���T�E��o�ɗ\�*�� Jᶃ��v���*�̡��>˃,
�>)jA�� c��%��tA�
����g��@O�A4����m��^�z�M����L
�1AИ��D�t�e���!
B+�����z%*����=eh�ɮE���rE!��8��&$�k�whCʻ��7J�7����IAh���lR�W�AD�е��>�!��~)��������9
;ĝ�2W�k޵$�A<�CҸRVQ<���x��$�} ]����"�E0�	bY��샭J��>{)g/N��0�g��I���"(�A~"_�ρY�T�>A�/��	�K�1�������||}=�|z}�,�S�L�|
�o_�����D��Y�[�zm$���a`6�]��wǭ3��6���;���"�}CW���U��=�S$����(��U�`A��r�a*��z ����Q؃e|�E#�I��0����AFt��J�U
� ȉi���IKe��'Xp���B=9��ϲ�����q���%t�pD	���!M�`ie�	������R��3>A����7�ğ������h����/6�0�ŷ�g���*:���M
�o���r~�jU:�x�����AH0�U��ō���MFG�{ݝ�^�g0���N�v	��W�q<�&�k��`P�V�	�����Щ+�z@�nhy�zM�-�_>�y��dc"Ab��]&rio:��U�S�এ	f]���B�� ����'�� 7�c!�P:�t� ���P&�Jw��(�J��7
A�4	B%v�T�Ɔxl��T�p��c5|�p�¸Ud3�ο�'�����#�O��q�#p�2H�7���!dN�@�� ��]@A,�)��3�u���	�B5�m
r�(||Q�H��|j�fq�������i�
���〟~0I����Vd��ebF�8�4����A��� _E�B(A�ELd�9~t�d�ie����}��y �&9iZ��T�a�2%�H��ҋo`x�n� �����sA�!n ��� ����@A(���@�/ҕ���FW�W�u��v��B����$ ��� 4�h���q?��/���
B���=�q'�q���� ��8'$��A���b����=;�Ф�D洜Gw(��a�� ��&�� �������\8��p L��o�F�ķ[s!gU�������E�1A�	���	�ܴ9{în�z	rOA?�qS�~s>n��N������Lj�BU�c>�'&�g �j�]�X��oR��u��/��(T��AN���|GY�<�+�-�"�XaiJrV�7�Gn�<�f�����C�Bl��}�,&@�N&�σ{A��vW-&�)���%��=�qVm@޵����A��>��PU}p0+��T�Y$�ZtB��2�ȹ�>���VÎb�Tq���w��a0;&��j`��C�ލU��{?6�Ch���U���������
�GO�C5N���4�dv��:�cI��)s�d�{�eZu�oЀ��m?�ۉ5���/�\ρ���]�OZ�\�L����=!�'�d!bv-�6/0<�8QA�VTb%ψ�@1+臼;Fݻ���^8�^�v��Pq���bB}�n�.<��L�e�L��,�ƽU)\���A�J�t�k���.��~����:��S8V^<h���&cQ�c[��L���Ą�y�^�j��s�� TG������6s;m� B[<{���J\x���N��,z���X��`��"�`j��[�FJ�#����N�Q8���r����"�'�腠3P�bK�&�,�uB�ڃ���d߀��G$.�u�b7p�{u3���1,��x����A�4k��'�����O�o<�����T˂f� o�F]�{�[�S�,�BTi��v��@PUm쎆�lA���܌����Ԅ���܇���Z:��q���3C4Ked�;ܕ=����7�
7/�Ql���ѥ����#��
�x�lɨ�M�glJH��!C<��U���!{�� T���	k�� ��B�p�{��)�2�ZV����6����F��Hɨ�x�6(!t������.s�/�hso0J�|������B�<����o�N�;*��o˗�ɗ���D� �!�m���D`�N
��Ʌ�.��O�Y� ��DV� ̴D�m	��� T���!�Oa�\�ހ�dp�W-�/p�����AԴ�X<ԃc�� Jfw�աyGm �ǔ̆���.������X<^��(<E��>�h��Ѷ�:Ԕv�`;n��
a�Ņ�@1�A�� D/9��	>���L"��� �ۂ|+�����3�&+�W-��];&�jUb��!LX��^�I��I��	_�t���'|��;I�(=q&*���� �l._俸��^�-^�jT F8^�	��:���#��!F%a\l7? �ō<0A��CnS�vc+Rj�|
�^��*C�"6dk�`��Jo!���
�'E@�LFtP1Y������mj�&�[�	���1��Lw%!���� �/�OA}���'a��s*�ś�P��@�EVwm�euK�L���E�Rx|�`W��� k���� Hx=�~*b��Ү�0�����+��|Ad��I>=|���O*�Z��]f2
���P�ò�/ِ��T7*ZBh���HA��E�aG��-ѐ"�r����S!R�ÒBC3�9;����&A���]�5uR�(�RJ�OQnn��&Bm�>������Q�����OI1����H�	�͌W���'�J���5�Г�������^ؔ�v�Ľ� ���٪dD�*�G-�P8\�q�V�|�����-O��ThE�� h=.��CnTUu#b�s�L�.��nzA^�MM�F��ԡ��������CBC.�&[⨀��T�XJ��h��b�y2�4%�:�RB�|2LPn!�,� ���$����RJ/N�
gR�a�%	�U�l� 8"���`�#���.��p@ٔ���BATB@���/��Od�l���~<�2��j�E��QX��P$z�� ����=AT�ĵ� hY5�v��׾X'BT�i��/�J�}C���{j=D�ZP�;Cm����q�p:xDA�wtG��� cĲ8L:�4N��[CH�K�1�A«�s����3��P[(�cD��F��-,�?�Ω�֐b�4�������� �?��	�������a�� �ډ�������&��K�/B��LP��:mb7w&���C�>�	�A߭Xn��ǻ@s>�����B� �tTAX�ȢyN�A�����2��7����[�W�%����ʳ�\i�^�=!�)0��
�np6�u+�̻#�Z�d޵�[A0��i <��
�"?;&�I�y���)Dv���wGଣ O"pw���靖�O;��h<o���I�l	�ph���$Ob�X������+��)~���!M
X�E�6��� k\I���%c��p�^J�x
1����Ȋ=��QZ�i?�!;��������X�������C^�f�0ʭ=7&�#�Iٽ')�ѯ�`���4���j?�&6�H�_r�l�v(�Yܦ���o��Gn��A)�~5>���ޏ>��!�9��ٽ?�-�=~��G���P���ϝr��G�Ji~��?X�wG�l��?$;�y��1~H7����cbA��?F�]F��ܼ� )H��{_����}�����9=����:��C�q���Lʢ~��?����K���P�#�H��a��]��o����H�0ʢ~h�>�;&?B�Zy-j����>���G�^�}��^ky}4Jj{����E�������G��^�|�����3)��3~����1��<���~Q�E�#�x-�G<0�ȥ��*=g���\�\�sI?��A���'�P{]�>>�_!J6�l���x-_�G�}V� ����~f&�M�m��|������]|=ȿ�����)��0�bb{}�?]�w���܀�?������@�SL������9�������ح��Bq�v���+��y'�+�x����Zm��T�'8���F�C�G��E�:��U?~�#�%�>�/��Z}�<���E�}W_.�ؗ�u�I��r6������t���.j�I��P���Mb�C���b��ဘ�(g�؄�؄��p�>~�����p9�9\J�����߇��E|��!5�������z�>���]o[7��ުkz}d$T��0��
�CnN�E���Y��Q�෎ϔu �����L]bߵ���t������=\�nO,���!�%��6�ߵ]uo�B�[�_����g�N�OB��j$����B��W�.���1�[�GT@�4.�͋��g�4l@�7��,��Z�a�|��yC7.rq����y3'��~������'1�r�U��:���'��I������8�-��y����L�gAs�ju6D1��ܓ�YH{��M�Me/������
�H�ݒ�w� R_�p�Գ�����& �K"bRd��6��Am��r��yŘ�
7�/"�� �=�Û6Xބ�έ!���Y�50�	�,]��l�z����+�P�E�:"�[G���ٴy%:��au���zI�s�w��u��ud:h�ݸ�=�E$';��A�#��ƒ��@r`;oQm�!�dN��h��"�WA�vP�v��@����R���p\eu.hxpA��1���&ڄ*Y��+=N��莏x����7!x"�J���+���u�
��o\ �ny�m�_d"נ'�Q�ѽu���0����!���E���2���d�^����9��09հ&{z�� э�-�P�T��6�#��1��mЄ	�����
�hA����4@H�o Ҩ��dsB��ھ�������92��L���ȁo�0Uyo�D�V;`�k�i���v���(<�or��Hf{�X � $�D:����� �H�)�%W�ـ �l=H��-����ew��`�
A��i����Wtd��y%ڀT��/"N�R�P	�6�9�0%^����( 	��ޡZP9��нC,�w�luJ2Ͽ��3-���w����$^Db�jꖩ*ϧ�:
��8G�b���W�NE>{ۏ7:���=�E�Q}���#�^��ɺ}B�O,���_D�F�-AW�D�����t��@�-D��Պ7�B]�Dz���C�J9/"� |6"���4o��wAX6|����7W�����S�8�^�~C��(<�q�������ɠ� u�;3�zlX� �� tm��������B�6�(A�m.�F���w��a�vېMZ�%� �ɥ<�L��<>��[?ԅ>��= �@��WԼC����z��@L'�f?N�ٹ ���ݟUuT� �D�F���-�oTZ��!L�AYsA��+� C�aM�@"QV�W�.@
S�Pt�"��#��M�@�8�*�R*m��
��QX������C�鋎 Ȭi��J��äo���k�=0�"fZ� *~&���VW�v��I�϶� �w�h��'%��OAOx$�������I]�	��RbB�4�9Z�7A���)���&��Ǥf���<k��-+�Q�����C���Y`�Q�T(��(46VwA莍M��\��Wq�:�Sű���qS6��4�^
�^Հ�<�9�O���t�".�F wz�� _}6M4���xK�D�1��F��ľV���#A� �M���M�Դ=�=�wՎÇ�� IjP*g>��z�;�\��P�S00���%{��BO@?�	(c�p�6��!�ħ �D���K$D]B*�5d��! �L�FiQ�v��(�E!������g��4;������F�A�=��@�o~&�#+e�9���PV�G��;���q`�7E�����q"R∀p�4��Y
ɀ��}�Γ9@�1�k.�Ҏ����=�����];��&s�=q�]Q��E����"i� ��I��ͫ��]38<Jh/R�oAx^> ��l��\�����?陓Ղ^֦�fwl�ȓN� ,MIĲ��^���[t������^�JD��	�FG��AA/�(�F�8�ℨ^P�5@�[ZbQ�qc�b}d�!� ���<q�X
�^|�n&��=��U� ބ	�3qL��A�P�=�<`!���&̙m�Bq�����9�Q](����,��GB�w� �M= TX\�EޠRt��F��F����� r���y���ZR�|F%��eu�����ݻc��D��������Z�7����|W��,�4�OF�����A���`�EZ�5A�$�}�[�[k��lMl���,�^�؟��X�Z�4^��kmEqA�c�Z �e��딺��J�7{���1�6n���T�CdWi��)(��M���Z��h��3����6��X��I� �X�Jpο1F!p�)�1qA(6'�n�Z�0��)E�f:T�� j�!@K�Vy��"%��:��k��%�ҡ�ypg�e����S)��E��C��g���K$. Aw�� �44Q����	��G���Pʡ5�
�S�j��1��]�n���
�2���i8���
���U;��Aަ�Ƽ��<��qy�ye�;�MJ�ɻ�Í��۾'T�:E��:m��T��@rq����V* ��U�㢬�(�Q��{h�Mܰl�>��Z�9@m�������Е�r����@��&$��S�$ބ�Z\��%��J$z�j��B���vu���C���m��lz0����B�"�M=�M�x0��rs�yUZLA�`ԶKxeђ��I;@(*��AhUA�C�s̝��e.��˯<r�<,WF�0��fdHn<5J����c�6e�C����@ ��^{A�z�+����7	QQt`A���Ƽ^b�%Aa�� �\� �P�T.z��H�S�KJ�a�>!�ԑ�%��HO�Nś�����a��1��-�k`s�5��b�/Nw��mE�%d�FB�gP�k q2���	��*#���s�ml��:D����$��b�0�qO4V�Z�ݻX���E5恅\�b�� tڢ�݂�:j�s��H��o�H2)�1��ƶ9�x��E�x��]���� /+H����ȋF�e�P	d��f��%�d��|�Aɶ�0%�s��I90hB����]���e%�����D^fP;6r� '��#����b��yK$�*��G$o��q��Q�7�i0������J��/"��Լk��AL� �s��ͅ=���� �>I#!ȭ\R�B4�j�<3bX� ?�I��%g��P�*� ���Ye�n8Լ�A���r��XJګڠB��P����l8p�vZ6kZ��A4�xf���Lz����`�w�A����[ZBu�7B� �!˯��Ӏ���Q�~��ˁ;iA����&�3�
 �?A(��9�D�~��64�	Y����Ԩ���F@����LM����c�f�B�*���D}6��
�Bc%y{�'Oj k%�l��=� �	ƀWZ��~�.-��-DZq>�5a`�ƄY`aS����3PB�Rp�% ����a���X�6ğr��))��ub��{R�칑6��(��<֌���]J^�&���S�o�nu3l_�t� ��f`�T��� �e�H?)n��S�Ҡ��!c5q���Љ���F)�� HJ��בpa5�`���y�*$I����(�rZ�қ"��x@�&Z�T?y6�ǃ��R�C�6�f�h&�r��\%���u�k��U�Cq�����@���X=� *Ձ@�f��\��ť �<b)Bq�"%��Rct�QO�a�8�އ镇���S��2&A�E��6 נ�*�am�^`�)����t�:w�S��s�v\�N��b�p�� H2�t���bYX���=a��I�{���6��QT޷�� ݌ |��a��x�/A|�%q��8��uU�%�Զ�|0V烑3��և��%��C�O���Ģ�=9t�&u���۷���ǧ��9�7w&���DR� ��E�υ袂��+��!jq-��³�y���]�.��7�i}7b�Ά'z6xO�������ƙ� ��q��o`�v�
�\@=��9MO �Hj��}��@�>��%.�O⠱ �WR%P�5�O�E}��Ơdּ��pyj-s����|�z�N�A �9��>_<Ԙ�%��%�h�ʝ���P�P����L;8������BA���hн������>ר��4j=�:^O��ש������C#�SתT��Q����z~h+=��mϢ&ֳ~|�Mb�j�?��v���}7�m�j磇��h?����`���`�#k�zdmR��]��F��lS9�,�r/~t�~h��~���kl���#F=��c����w;�?I�,����}7��-�}bg>zxk��\�������͛��cq.�͹?�e�W�m0ڃyCr>�]�'�����烱?�✮tX`��ݥ1�`?���R������c��J�?4׏6������:��q����{q��f��YVJw ۼ������s��?�b76₻���{�U�G��`|��C�M[���<7o�S�&�����R���t��.�#uwT/���4��]�D�~*SZ>�t�I�5~h�啋���%��s�ϻ�x����{H���B��<�bm;��ݜ��C�ǰiz?T���|.��w|NV�ܛ��B�[�?)�׀��ҽ��
Յ����{�����f�r � NYC��۔2�!��S�e1�C����Bg�f��	�=.�����i�G���t9 �Nf���&��^�x\h4H��Rl�#�����Ͻ�����M���!�q�"f#\Zg��@��}�����͙�K�}s/��lw�"�t됏�^CYU/yx�LH{͉����{=s/9\TM^�?s����1�:�ٺϦ5}ƭ��hk�LY�s��Zדy��\�mC�rC~p��1��]zqCrJk�q�e�v���>>��z����h>O���St�������n{c෦ϋH�
�s�mT�؎qA�
�2d�<���#!Å�2}�$��΍��C�ۖ�]>�t�Q�C��p.G�������^�/�3�b�D' A�_J{��$h�B�\����#��t�P<��J e��	��̓���P,�AL� ��d�֐O�J'�!��0ѷ����@?��V�!d�j�� �C��l��4���☫st����ǂ ��]!H�tP��<K_~�+��^�h���xPf������D�>��`�k�
J)�%B�q�W�w����FzH����q5���H(�U|�C�͆fӀ�� G�!N�٠i8�o!s{.X�	����SY5
*�^cec�t[��[ �oW�mE�8
�KΰÂ��6�rچbKiI�go�2���i���/��A���=z�M(�k�7� �k���u(@u�*+%�S!�M&�$�~ْf(;Lm"�[_DPK�x�� 
�%-����j"��{PU��JX�B>���:t�.�v����`�F��!H�<����82Av�Q��!�����!�34\�vJ��N9�> ��)zC��ީ��'ԅ:"@:��*̛�S!b��,�A��rA��E6Oh8D� �s�O�	)�>�/�w}����X� ��f�:��T�J�����D?��]�`�,$Y�Y�7!S�B�fa�S��B�t�yooҖ��C��3� ��e\�C�0r����#� ߝ�z��D_AP����@�ArZݽ^1}����!*�h�����7&\2A� ���I��?ԅ�����ɞ졄�n��^�'�y u:���N�3¨ /�t������ur��0!��L������%ng(�xD���Y���X�gS��"O�٘'�����R��7�	�i5x�RWn^�?g��D�8V��`��Xz�Q�w�C�"�uو�@_3:�
���ڗ<�C�P�@D�Ջ,9o���0��y%��9H}6�"?F�5��.M���٘8��]�ЄV�`���X��D��|-�~=P=Z
$�ca�:�p׿�*�%���)��p0;Nj��3�"?6N�Fd��H��kC�`ld�i�����	�)p�9H�>H�.Ϛ/���ښ�0a��7s�0E�Ǒp�A.!m/#:��)&)_�mI���HZ��^� r	ZÂ�^T*Jl�� ���_�����A��`b� �h�ԇ���m�Ӣ`~/u!����i�Ft>t�k���O�b�9��oT��r:��n�l�I�F-�v���T�lҨ	� �(���&�%� �°� J�A�8y�1���-�����r�"Y��P�AY���YT|&v��61)y17�S&����/-
���%��4���"`�'N��`6�~<��&}���"�q%U682ը�.�ï��XABk/��h@�xv� �⣢�E%�=7\~A��H�.�+���e!�W,
� �j�?(�<x���TZ����I��M�	�
�ݏ6gN��fB)R.��+�  ��H�����	ʬy��U̷p^8+��!�đI��,�;���A�� �s��E�(<X������e
!#�P��1"���g�?C=V%� H^4,ړ��Ր�sA��o�͐ he4�3�����TB�&kA^V�8C�|��'[�#�gu���A�R��T�8�Y�H����I�A�Y�k����U�C��kR@���B�n	�ʤRѤ�Ǥ,9X�¹\~zw��A/������X`�X�jL��Z�xl2����L��g�p�J$��v'��0� �)ٳU�����ݠ5\�s|*�: L��r��+�^r6>
$�+L��:V}�+��)�J2`���H�c�*�d ʻȅ����k8V�%T�B� k�x�U��/ �Z*��G��p���4��mA��M�D�-r����RA����!S�2���|Z�j(�� �D�A�'!��(���� o� �(�GT����Z0�а��-���0��1�4H�~	��B��)iW�f�������A ��Cq8�� A�`An�����~��p�큃�M>�=�!.Zq��@"d� YĞ&�A7����q��yCOp�	�*��Q��@S�UP/*WL�+�R�4�\5Z����{�kK���^���ԍ{!zM�	L�2�����@o��ͦ���MR���o0�SA ����9�7��
B������+B�b)���q��#��M��Ү�J��ȝĚ��>�N�R%����Z�v"��H�=� �B�&>|O��Y��x�������� h/l~J@���l<��v��J���q��� �� (<�7eA���u��O���a���
WY��MX��A´ �ns��S�ַ[���@=A��+d��� m�̄�����;�$�Q�M�P
�� ɠ�����١�0��`4im2�%&��A����A,e"ܠ���bPgC��� j�y�n�X؋j#�_\8{�o��	�p
��f��~0��^���"?O�v��}�odx����AP�>S�#�T��1���Cr,n��D\\Fp�."��$��� u���%_RfG�k/�S%!�(:8.���Sr��	���x�.tp4dȋg^E\��sp����8�"�'?��8Ha';�^m��$$@u�|�|����X*�B�xp.��W���)�fC�� pn7Ē%�K��?�uc4�D�b%H�_ɔQ��!�*�>K�߈UA��/A����� �˸��~<��Xr��\ё�]�px.FvD�f_�,����A�qțj��q_��P��)9(8$�*+$B���c@e@:)�X���8��%��lOsR�F6�%�;s��B�Nf	�s�A�1�ģ\���S����V]�;�6F�
����!\i���Ȅ�S8�8�����Cn#�K:�GgЮ���Sh�,��(%��<$(W�1<|)�	���րC�$R
B�9K�*d�����x�_wT�݀>��D�噘|���@� o��ȮR��B��4�>Hv��|�O��Dш ?�C��w`���A(�����SJ�?�A�����4\[�N;���l�E����
���;nOO'�{ǈ.�/�c�*\��������6�}�/��'<njπ{d���c�C�A�4ʽ��C�R����fYM>ao�� �XAn����שc��@VR	(+��� ЃO�ߗT^Lp�/Ⱦ�|\�}/Ou�~�2[&_�9���ʮ�o\;?`����et讜��T����L�X�Ϧ��N���}�A������R/>�|�Ց� �je���!,ҥx��J��$��j]ŋ��<I�AP<�ɖ�h��0��$6�'qt~�"A	��b�� ��Ρ�K	��@�e:��>���P� �@S���\ҡ����h���CB���A�U��?DHl�\m��k?����w�������w�{H��֯�˕A?��v��H^�&	�۽��`$%o7��������$I|K���\,/)��/��ȟ�&h}	���HF�Ѧ�ĪFQ��CH�߽�c;|��?����WE�Q@ H���p���~al�1H�?~����<������M�7����}0����3�p�
��3Ц�h�'�+R������_�(Ü��y��>b�[lӹI�?���Õ��8�!�Oۇ���\}���T�!�y����}S��b@�^�e(s����^����_㝍��{��}}����35�6~�h&�E��������&+�m����~]��KY�:���C�a�C�o-�z��%��?��{������r#|>�&�����ݿ����Gq	����_��R��+�G���i���d���x����p�����g�n���۝1���6�,���Њy�l_��nw��gR��ٖ{_�r>G)/�z�,�˙�{8�gy}��g���'~�8�� ����j/2����g^g���#��#��{\���U��y6/g^g���U���r&��s����鈷ؼWmH�.�<�߽�s�H[^$�>���-�&���s���}��[uW/؏�y��}7�j�{���l������e��q����UM����Ng�߉g��N�5>.����wN�+��">Zbt�Ҙ�bq3^�-m@����"�b�$�{'���7��Ρ�	��C0�s���.��?R�6�����U��\W-�G¹���+I�4��
����>��xۑ��,�p㷶�a����zA���9��p��B�yµ��?n�r�]m2�h@��T���$�w����P��/ oL��?��pǂ����B�P��(|N��Cm�1tk��k��r�1)$F���C�z�� �ZǱ}�8Wo�c�M��U� �*�ZG~CE�{w���~Џ��Į�[A  �P�h�Cjc�x�aʿ�CtA������y$�<"�<j����자�N��ep�Oʶ�o���(� ���I����z�	¥��N/�94�����N"�6��gTg>r���}Q&`�#���-<75F�W`�O�EV��A�@z� ����x���;^���v@2�y���O-hbP_`x�� hꖊ��z1f\&_$u�vD�&��	��A�''�D"T��/@H -ah$Tg���i��w��<Z������v@��8U"��d���'��pF�F��	���X���jT4�>�K�t�fGA(k�`���PX�ĺt&�wu��F�Q������AL��9����^��-(��~A2��J�g7��7�rս"t" S�G���I�BwzGĨ JZP���+�w6a��N���!A`=���(e
������C��%����� ^ZaP�@$X��W;��غե��� ��O�	L�q
��+yO�9�8?���)X%�_������ ��7;	/��` ̄��)$]�Q��<A0V�A��b����_�#�e��)��F&G�����o�u
i���M/���as6x{p"G�~�Au&:�>��у�\n'*11������!%���Q|B�"� 6'@�U�A��O$����eJ���Dc0%�}�|�'������<���(��P?T[:`b�U=H�-n�U�P�o���|�,<���ʌ�bF��-���QO���Epє����[Ax�L�g ��m9!�o�`C��[���aU(e�>��% �jÑ�h�|��
�:�n;�#WA��P�Q�Cd��а�!'kE	��'H�KvDG������<��A�d��T�/�cpLhA��l�(I�&��]29���Cr`"�V�ܜ�� Ǆ[P����v��ʠ�����0[A�	�%@]h�,�����/n�Bl�U�l�� L,�� 1�A�:������;�#:�Z��֋j^����^�r��jCb�]��x�H#qI��C'�F�f�j%��Ի���k>pt����fQ��������������r@CT�l8Ĳ0��I#�/B\M��� �E����)��úO^�^�>@����Q�Lx
ۚ�a'J�O%x��wBs�ns�TQg F��(jiaxw�"����a2I��ʂ٬�  ��3���sr��p�\��mMc4�<�r�Ԁ��X&��\�h��X �\~AdQOfaC,�w�zs27n.0�B.(�j���-$��A�ʆs#� o�:���"������&�:(B9����/p�8,��"�ߘ:7	�뒎��0� ���y�	j;��s��e=X��ٖ(�@�&ȷH� �~5'p���ʟ�J4~PE� �&\)͋�"9v��]>�F��(f4\��Z����w�EB�Ř��qz'L����}R:���//���y�%��M8(M2�0�*j=���5p�+u�Q�������*���ș�<_Z��������&uW	9�#�Zs�����E�p���	u5���F����FD��x��vm0�	�m&�A���`� ���P����kC�y�.`q�+�:h'�c�|�Y�ʂ�Wu6 `'ub��'��������%��b'cB��'A!���I�tO��E�J�	8`3^^�:T�9�MZ*��%
�$��уh���଼N<�PU����Lr�y�~6��h�-���Rmp��㵂��_AP�hߤT.��o�dl
j�?=��}j@��p�&Mء:#"!ӛ���F��.A���g�7�0����Fi� ��������e	a�гC8������{�+w�g��O0�����C*6}�=�R��#j?9�'�Q`;�r��������b�ŉ�����a���a�{�dkoJ�I#��M�����;6�tdU�C�� �/ @�����`��$K�P>	���dC�Ig��C�m�zvA(B�;��"��aB�T���}h������A	fx�����aD���1���ju80���� ?Ј�C�#�x(��Tʡ�3?�g�T�j�������T�����`�D��DõX4\�	Bw4DZ����W��iA�N��� ���
�@�O0�I�(�xw��F'��v>�D�NIGx?�7��H����w��(� �I��6?1��� ɏ�`��EILPu	�����fL��8슉����(���5h!Ϊv��A;�X��,�C�-��U�x �`�8��%���q#�*x�ra���`"b�"peT�מD���"p4P��>����b�*&�["���-� �P �+�P�qC��&Ɇ���#!�Xr(J���Z%rO� ++�W� �KF��'�P�*Ώz!-�ǝS>�x&An��RATG �����"��+�|ۙN���L�y�"�7���
 �+����g�%O�7���^�WQ˗��Bw�-R�NB�N���p�B�����z���%L  �j�Ǘ�"��a2��-@A�E0��|o��݅0�Ʀ�����I���Ƥ�UNܝ�[���x
%E��-�pʟI��暾����vA�����\�~\�	,Eo��En��&6Q� ���������{�z!�:��+cB�<!�
�N����30�%[A�	�7�����W��qw6x�$����`Umj��p0
_�Y�oA�$�g�@O��\�#�S�0�AP&�wxeT�>�=�:3q�QB���/j ��*ݿ�lT� �\�<�Dd�.�<8r��'K�gE!0\��D},s��O�4�h����i�X��@�������u�i�L@%`s�6�������wH��������}&A�4�Q�P Sy������|_~O_�aLt���#�C�&A��%; /�-ҡg�M�t�3p�+�e�����x���S���B	9�E0��I��0�'6ć�9u/��8qcpI����E��E�xAx)k%��-��:�&�!��ȂP�a� 4ᢲ�F�� ��AK��qcK)f{7�D@R��U$��qUz6
��C�T�Ҝ�xL��U�0'�$��X%״�jt��G�-BX�;�
Lŋ6:�V���ړp�Qs�@(��O�1�)�������:?hʟ�\B#M�sT>��A�����|0ҙ?�Gy��s��w\��/�w����H/����Cj���W��6H��&���=r��4P.�T@�g3����m��P�`��.������v~I-��?���{�&]}�?$~�o�2O�w�燤�������|�_�1~|�ؔ���rJѦ#(1~}o��d8�Z��?��1>�y>�J���|e�uڈ9(;2����1>�f����?$K��2�`?��g�tÇ,�Ѿ|�>����}���A�����_ɀ��?��+����K��I���~}���Yd�מ�:��*}�� %���Wma����ȆMw%�?_��`(֘r	���?!���[?T!Ρ&E����0�I�ss&?���#��)1�8�U���+�H�?I�c�z}�?��w0�@�W��B��N��.�8rY{;N|�ч�#�\��?N���=�+# ����|e�r�@᳸��W����d�=�D���������d�5�WX��[7t�JXH�?�^/a��������A�׏ӊ��i��C��0� �7��,p!�J�5d9��N�>�S��py��O�����".����+>��k9=���]�G��
H��B��ӬO7�A�����J�!��H��n�p����G�g��C���+�v�L���H:��#qÚ_a�τ�!d�o����g�����w2�\au�������"�y~D�/b#��҃�#/"�qx �qn��%��3n�����R! ?����> u)7�	Y,�=���r#OUkH�z����ߐ,�� �l�mZ��{�y{?Z�/t��<���1փ�}��_9��Voh�}"أ�@U�)�
�#��i-��'m�C�,�t/kn���)x"�Qn'�va`G�_q� j$,�mZ#R[d���X|�x(3������8�X������`��o�$m#U[�C��Wuo�����T��Bz�l�dh����1��AU&�~�mB�B#�a��<�c����Q���=�1q�TB�ު���zP{&��P��:��x�����$$D���GC�T*���F�W�|�lp�rM��'@C���ضAN��º��a`� �Z-��u)sn(
�:�z�f���$�(����7����3��wHM���Y����hlՑ�>FdT'˃ P�N�+����N�>�x#�T��*�f0Q#+���AW���Er}f,v���&A,���YM������R�)�a`����#g#��o���0������,�A�xP|%,�A܌��1�_s�#|��X�2�^�uU����XW�:��L��U��]1(��Gw&���\1Ah��h�~صg�/W~Q0�V�É|0���`�}�/���a<�<ُ�Hҋ�O�����eMpU2l���Hj6�� �J �Q(`�3��kO�#A`��|�,�|1,v_��"�m��[]A���*?c��?גb�����c J�ZO��'�4�v;8Z�:�ۜ1{;&"y*G]�x0Z�	���b!([����n���a�/�?(�����/�j��0�W��wP�@Xt7���|o���È"��z"N�G��Sla N�x��0
�%��� ���N$(�9���ۛ��NY�����-亭=9�����Y0g��ga99&�Z~Q/0�	C��l��H{�?�
#r�eډ�C�AV�6'��m����l�u���E�d�̂^<�O�j�R�t��Af4��??J�enG����qv�+.�?h �K~q�te�B���V�3����#�~!p�r_kw�6��75!	��vbo�e��qⓂD��O>'T'u0k��/2'���J�$�d����cbc#5��������6Z01�6�@f@���JA�߷N��b�w��s�g�?�h�P��f[_"o� ��"i� �}&(��j�@M���۠n@�A5A_�� t�!g� T�Ĕ��c1C}1�j=ȷ
�g��*�����׃1!��iG2�*l�W��pe�V��������I��
�0��:��.n���0��(E8�;���qS�:��;v��t� ��C�]z�Corux0��k� �\v�*�N��f����1�&�6�^�:�5 Y�/��Ֆ�2�Cv_�9��:!lP| +�૞$w�)GY8�.��Ġ���4ja���|հD��(�cu-J/P��{��l���`L,(e��)#-&`�M;���>E}�vCj1J:m��hmܺ�<���n����E�
�ֵʂ�
��
�r 1� ������a:5�����$�sV���J��ɩ%�2��%�5�L�w��,��������:�A��b��d�u +��� J�¹x��Ը��$�
X���)�M�ݰ���v��k3�[���4��I�����qҼ;T�7�e�E��������N�f4�8�ħ��ڊT�S���w岴`�$��ֺڎ_�$w�~̷ۍ{�܂�j�0;V%�b�.�Z/\�l��ު�{��r/���x��TWAO|�-�޸O���u�U�Ma����Z2���;p�$& '`^ہ\}����ّ�v.�	S�n'���֛0�S�q�S�?U<u��3�~pи��Qu�``(�Z������{��&E:�V�`PU<���Š��@�%��jBVP~G�`����X��DCVy]֠x��q��H-Y��莎 fAnD��œѲ��"�vkNM�̷Qu���I�8�/��@�8�����1 ����~�5������X��!1IL9!�<Ȏ	*�୮ V7�A�X���r5t�绪�nA,0����|����T���� ���x&A�E�f�����(��AA�"L�/�n=��S0ۂ�%�ݍceA�h�	c�A�_����w�P����@[4���VMP�F"a��bA�A��$�r��&(����~Lr�&ؓ��	B�Hl�#q�.�Y�В��@�3��]S0���q�cQ����%5-��>��AGN����pD�QY�7��#Q,�D6�xi\� �َk���&ٿ��G�Iuwy�~4 ������>S�6��~�����Bp/N\�־ ���-.T���v@�ǝ�,�B�6�C O�9��SGi��{t���`�m�6: ��`%K���CvA`_� |��r����Xn-�7!�����VT��K.���Md��9���:�DH~Qh�Cs�ȓl��ˍL\[�.�����$�yJ�%5Q4�a���P��!{������P��� �v�O8!��S^L�2�G[X��iˇ����l����S�"�0��;��`��t���0��7ק����)Ar���3Kv�5��8�5pmqz US�go$�ɱ�U�4!r|t\\�ބ�.��3��^*NH�Ib�s�B�r�
0̮�����oC��l��X���s����+6�/)�ʬ '$	l7n2N@HP�yI&'H:p�e|��ڌ�E\���� �o�tVh"�z�H�7&.���t�Hm�j�hA�c�=_qBb%����U���7h`i�7ι�����/��?��6��.�g�Y?�9�kg����:���,Q��ȩ�.{���Gy����kH��v(/�ߥ*�Xg��N����.}L�n��]_^C�ƕ>���~w1�X�(/p^g�b#�M�G�� �	F���&�����<�������=��`?��t��~���Zg��wo�>��?���j&��̃�|�)>�`5r��N꿢N��h���v#�\������J'?��Z��z]�J=�:���nB�F�a�����C������<{O\3�Y�GK1����s�$��Ly��,��d��I6�6�6�K'��q3#n�z��gl7����v�����{����ת�������G��..�S����"Ǒ�Ʃ�!���"^�tb��p�rE^_T� �k jk�ɸ��{	�K?�//a�ST���}�>i�K��H����"�>��ظ��r�_��F8��'������;-��N�5��3A�8A�5��%��֘��r��N�w�Tp=N��QRz��o�ڋ4<�g�ϔ>~�e_y���}׾Z�/��NG|<oPb��{o���HB���'����۽��{����"^�>�c��{�"Nw�~>~���:g�L�&fnn'5��)��E���L���d�<n>q3/՞��5>��2�JL�+�0�T���/=�#�>�CȨ/6h�=z�#�,}�/i�|��ѐ��
�@���7QU�
�+�֐���Ƭ�P�y�L���)2�!۩5D��$$��������ؐ�,��pbTΈ�#��*
����h�WW����_f�ZG�_�PT�_��(fE�F9�D(_Q�)��*��;Ah����ob����يj��_!�]J�t���*�p�("y� �~�'�OشK��<~�V�g�D�|���$�~��\[H�nT�n	v�c�$�A��� �!�ZZf��pZ<���5Ec�I�o�EH�@�i$��@�P�>�8��f- �(Xv�����R�a�WK������t0V,��MQ�xHk7�6�6^�
��8�zș�����-�Y<��D�� ����D����<����y���D�q�?�A��Q�ņ�����S��:|A�E��!����L_�C�u$AħеU> 0�u��>�^���O�z�I�@���y!�3TM���QN�����c�D����$`1����0
���H70��p����,WEg���	�3A��$D�������]`c)Ԋ�����Re�5~_H (����x+��!l�䥣�7�J�� 3B0��)= ����Џ\���a��B�x� =@�R�J�v�6��t������3�Hfm"��'���iK�&��{�-P�z�{�xo灧p� | ���� ��"t@E����ċ��f�I�rP�ia'�Ӽk���y������ (h<�O�5����Ђ��ذ��*���R�K���$H&a�GG�����h	b�m��;:��Ò&�:Y�Mۂ����� &(��x��`8��v��$Zc��x� '#H�Uw�	�sL�FM���r[�A�1a��"��B,TQ�xK,�dV  �����4K�Đ�WϢ%�p�|llE�� �`�D*J�np�	B?nD��B���刐�ģ�,�8�+X0]���f�wGLw���	��H�4�G Ԫ�P��o�S6Iޛb�A<�?	֓�`qA��9.�M���#-A��5�a�`�=8��� s�88K{>A���� �a��R�H��m�P�1�\rgw{`����
U"E&��N�g�n���"����ų��x��l~ԅ_���/���$�v\�,��!j`�K���C~]�D���� Q�.z�K(ov�Zq���_�N\3�s�Ҹ��_��/��pl�������pG�9F�V2b�Ƹ���r�!r����ޱ�7��ޚ��<:��|��L5�ׁ�L���iq?�rb�8��_�=��:��3��r�o{�;���� �e���W��9xЋ*�-"i���'FN=f+�f�����ױ�w�ǀ�'��Eo�y����	q��L/�G�ӟBc��Q�N��їٴ�*�/�,L��7t�^������n��G�|���]N�BT2�l��O��`sV�^�޸l��A5
J�Qز�<�Q���52V�8���bq4T�A$���������n>�37�����躲v���1N���Q�N�ft];Z��x����1pS�fR�&R�H@���Ic������O��p�����'�>c2�s���B�����p5��B�"��Y��;2n>u�׀��3��S]�[o�����ri)��f��땀��I]ȣp�-/���#?dcc�2�K�r�C���7�u,�U�K��:�x\�����@�9b� ����mĦ���O����z��Ȝ�0��*|���8�J������w��<�o�l�w�W�9z���������֊�9��w�ƚx���-���װ�����˘���u������ٰ('S�r
�c��BzE��}	��ǜ??�N���_�H<ணd���~@y�k�D��-zLK����?�C\oN�f���pH���/���[sb�6'�Nsb�~Iu��M�$�"�����0���t��Jy�++�~a�?7�DS-�B<�����,- ���Q��dZ��97��K�V>��F��<�r�H\K�)��ge�Q@ys��Lu���^v�K0�l��=P!�l��(��cR��\y�Ƿ
ı��7���X&���d���$ ���	e@�fV���[K�V%�rU�=�n��T1�į��羬�^�H|'}�1g樉�\�X����f��`����X��j;!Q�w^m'#huvVG��cyG��l���M�y�=Z�1נ�s�Y�X�s.��נ��y1�c��=����֒�q≽&��5�y��,!:���7�ԥ���km-6���H��E�hm���r[�F<,7T��al�ۖ�~��p[������:,�'��B�K������Tq�����=���ŕ_Ƕ������]�t(��]XH��*ol\ΞP^��Y!5f6#v!�g���� �]�/�n��B@��Y�(/�������N�"���|�fo�Ȼ��m��\�������n7�c��K���)����[�+�ı�54�w;d�a������]������$�"�"�<U�^��G���M�ߓ �=�
�d=m��B��2ؓ�����霬��D����J.6�U�B}�|�,�_4��3��|���/�>�������fRsM&s3ٺyn����}tx=�-�pO��s��Vԯ����B�}롈PX��;1`��]a��.t:��l����/*�;�2�w����/d�Ś?�Հ�p��u��f@����1e�yU=�����}̵���ȁ���FQ/ ��Z�짱�s$�e��C��:�Wň�#���h_���_g��tj`��C��s�``��@�1����0�:c��ۖ|��3mrSS���R7 |'!���γsb�:�֜����Iu��:�Yvi���[ga�7�2�SjE��颴|�����wL�ȿ�) �fB��F�{��N6�����T��H�m�s(�_+J�)���m_�V ��9�>����h/�C[��}~L,����|K���e��?�)_ϗ��%�-�����b������Y���k��ߘ�ǻQ�1�����|0M��Q�xGuhZ�f����<s�a�y|~������Ĳh4��|����
	���X��O�������b�������7��&�������|6w?��o����_�yC�ޅ���卦|��U7�~��ջ}�,_۱���;��}�'�{���{���y���x�Ϙ�[��r| �m�����},����8��ۿx�1�֞rt_G|��֥�h��Ac�ΞY?)�_'�?L<���yȯ��Ӗ�y��:߲�罿����@�?7ʗ��0�|�O^��������_yq��o�����z�lLYA����Y> =�jdʲ�=b��lC������z-\bbX_��ϼ2��UL��E���_�.���rd$_s{6?�l1y��	�Z�a$�^��?dc����`��T��63�M�(!5[�}�?�KL0Ǔ�<���[B�"��l��O6lO�t�d�H6�|mw�!���3?�1����+3_�؟Q��v�����q��Yg�6?_��?�򫷤���L����N�a���/���׃�e�m~�l��0	�����5�y��r��
?$�-1������o�YBJ�vͶ���`��m��=����g�����r[�;���x	��M����y��9|_����Cz~�;�M��X���z��f���6��a�Yq�|(ŕg�5����=�`��X3��4��wP^��ұ�+lQ����@p!N�5�Ħ�$�E~Q@��U|=���R�@�J���("�T�@��B�+���x�X6[��x�f5�dO�|̰_�ٮcm�d���N�k@4�^�:	s��q��ud����WF��rt^c�ˏp�iW�.cc�;�h���b��߄.�*�ȗi#�5k�ʄkYbU�_�۞o��x�B��n�!Hae��{29���V���p_�5�|�)����P�];LNǥl���{�Dg���k�!�a�i&G!>H�M$�T� * ���ħ���O���ء�T�/�����a��4<�
12�z}�v�o\����U�,�Eע������̣g��Z��S+p�g���q�ZBayp
l8�)��0 ���]�Z2�v_�>t)��tp���}��[;�D�B�vj�O�D'���o�������gb�3��HȪz�*�6 |���a'7��LN�^..��^�5�,<���ą* ����V�=�9h���m��J�*	��oX��qۋiT̆��.�(�.�����T]��K2���Bƀ���ZE��A��лn`uCܭ�]�ֱvc`���op]�QDSR+��������|�D���g��|�AU�&n�S��AL�bP�k���Qd�h�����kك���"b�@�B8>b}��05�d�*t��aɈ���M��ƍ�����1�m��ͧop��Q\�K��p�jm��켎ά� j}��:�;���Yn5�5Wfĥ�̘�s��m�`Ni�oh�cD�5\����4BLj����`�9�h�@է1����5ߍ�,��������Vs�W˅�Js]sS<_z��ভE�����u��|V[ȍ�m���u0?���6[)�T>�S1�TW���Ms�f�n�U����N�Z�垩��^P���*�J�����G�ݖ���M�^�ܯ�?\�7��<Cx_�
nuZ�`�Qh��^���]ac�7D27v��s��\*�{�O����fu�ѽSD��w@5`a�6�D��D��w{bH��vWyҕ����������*^�=~�nT�z9�'w0]�G_�Xt1d�EbS7_������X�9]u	
H3�F[�eM�Ǎ��B�Ml���{�h��&E�kf;F���.�5Vi�������h��0UO̓�0w�䲡��R��<s�����b{T��J凅R�]cM�}T�x����q��2��thp��\�Q�O\(?�J3��z�ID��/���2�hw-������f��aQo��Q�]��۹����u��7�qA���>{��G�V\�Ƭl<�������ք#ųK��q�<���V�!6����5���aM7Qy�����	) l:�䳚��q#2t��ݨ��Q\�<\�\��pg��Ʊt_[�.m1ňu�nu�?���N��y���A�4�6��M6j����<�K���a�v�����8��Ǳ�p�.�8�@K���=^��l㣩N|/@=|0���~�����|�����:j�|���,�+�B��Z��CB�.]/ߐ����T9�D���zy�B����f՘�Rɘ��4�m��r!NO4�4O6f�z�5�����]4m��Sƍ��(��Y��0�k�]O�X㏧�Z��uF�q��ǎK$�P�͎��8��1�qT�tq��o��)� ��b<'��as�q���"�% Z���4 M���W��0�����\,k��]���h������`��O�<�hJy=4ۤ�P��:���r�VG�<��D�;�خ������*(O��'��]]m4q,�&"����tN_E/�B(w�ׂ9��x�ųu	`"Am��U��{!��Z�*FK�K�U	_\M*�q��fxM���( ����aذ�ȣ�u��/.�ʴˉe'�x�������_�����q��x�14ym�O������X��h�����j�sF�yz�����5�mDc��Z,��{{x��`�7u9�Y�vry���G�]��5�F�)0�#�gM2c��g��G1�]%I>J7�kM�w��˹�n���F�\�.���!=8 ��~񴣜�!�tN:��b͗-�\��+b���0����Q�������w6�v�����V�Q�:.���ˀ���S�kM����:���z�o�i����t�mwt�{�V���3�J:b@���%�nM�9���j��p���5^{�m@�qӿ��p:����::�ٻ�3]�n��h�hӲ���cC�A�g����5���NL�d��5?��1��[������������\~C��^Ȁ.��_�"W`/� {��z!�bI�e����>'FL ��m<�5 �Ol�<7����x=�p��s?�������Q�y&H������s?�d�#<l ���@8����}�8&f^bj�z}�9�8�i�W�\O;��F�q����t�`��S}��ƴ��'a2^6J����X�P�U����F��B��as�s��k�/�4D9G���nDS��z�_:�ҷ/��Š�:�B��K�`	~,1�<	������\�����Qù&R���U����铘��l|�7��=}��_�	=��<�Cr��`���3I���x�Cܳ�Y�Uir��
�`%�{��iN�� =�Z���;n���U@@�s?r\@�z�l�*�=����
�0���CNH�>��^8����d�-���M��NE>�rZ�}�?^����y�w}�����M��`Z��w��k9���6ys���]�Vc��Z�b�gU�{��ԗ~���\��t��\߽�ז���}��}|����m����_���+�bM���|���}m������Ws��~+���h�8��xG��m�&k�o=��x����b���r?i���SVv�h�|��?Na���{��H��y��[}޹��S�������z��@�U��q�i�����[{��3!{WE��_������ҲOOi8�����o,S��1SKv�=���7b�r�;���u�[���?d�k$������&���e�-����>W"�������Og��	˾e?��SW���׫';ƍ���CVFp�m���ļ���~���s����\me$;-��+��r��r�>[�1�o0��s�ɿz���[=]��ٷl�|��)�����V����}�9le�5���z��?ϭ|��X2Ռ�缟�i�+�U?��[�ƫo〸�N�:u�_}���!#�����N1�"2�z�fo�G����3�(���qv	y�\(�q<�G㣀0��~R
ـ�Z�X�0�GQ�[
����w_*���fc�-�ZKe�TD>��R.4�<�b5#���I-�����ba|�R�A�]@y�Z:$�+���	���h�}�0u�r秘P�imy1)�6�ˀkuä�
��(��`+������忢(����'1	D��P�PQ�yU�~��r��,XA��/ޒ NNҹ�F�`��M�h@<�MzM�(8����IK�CbC�.���r7 3�񍸮�"�$ �ح�u��p�yt�y�=�����J!��B���	C���IaG�]{����i�$
��z���2#�V�19��p_�~�$*�k�����R�0�Bn�!-���NU[�ڐ�ݡV�%\�z��v&�S���WM��z�(�p���a�.���Ub6.+_%�ʯ�Cd��K�ϐ�i���z��Y'����@P��Do���d
[��k����u9"﫮A/�_��ـ�6���<Jˬ=�7\��~Uk�7�1�І,|��t&�����o�T��Щ�3��:������t�OG��ܡ�֞'�Wۃ��=5�;�CvkS��� W���9�Wƒ/�l�
�aC����������9J�V�yU��8�K��Y]�!~�0Q�.�ΐMuP@yК�JM*�%�'�+���s�(�W{�u��&��B�0��7�K#�2n�_"�x:���q%�f8 ��>�b�3o{�P&�7k�m�L��מ���|�Q0�<�_K#��pik��k��N�p��{}�����/8:m�:׌9��~b�q����49��j7��Xu���Q7^a<?�j��Na��;5�@`���{�A�p���|Е�@(~�yg��߀�D��h�s�u�(ϐ��~�����4y�+�VP@�����hV���
���3��8�B�+�lBR=2z/���O��Tir����q�L�o�u��XR�g�u\s' �i��z�Gj�i�V�q�C&\��}��T;{C�9f�X�'L�Ѧ/�kci���s�`����5���>�`�C��������U��%oY�I|W
ԧ�G���>�'��GF}1��K3�+��vL�r��j����or���l�=�G��W�u��H,�^^�ʓ�~`���6i?��F�x�r���l��0]	��g�g�K�HolT�)l��S�7���(�u�gG�^�@jU�M�ϫb�0j�=�\�(�RF�`�j�S!N��fp@8��
,�c��0>��>����u9�_���}��&�n/��1 }_sUl�J�1�̓s��|B"�A�Ѭh�|'�⇰-���͞�J�XHe��<l�������+�p�$0��+���i�q�hZᾴ7muc3�e���a.�e��Ù7Sc���8(����՝����aKq�iB�6�����*e�:�g�n��B�E@��]�|6��jQ�gY8���~rYJJ��S�����Pa_(O�;�[O�2���O���a���O��g�z�.�1��	nBYw@��t���%(Wԧ:�iz����Lx���7�ӫP��O̬q�D���� 4q	��>��М��o�D_s!sм�I�k:M��c��k��P@��S�cr�\HR�fG��0�a! ����Ƙ�B�'5sO8��b.������y�l���e3\?����V�����;�&<KF3�4\{X��Í��Pš�*r�&�rˉ֋��n	�]�%�g���d[���ѵ��o=�;^��6DX��V!�o��;���}6
<������K�Ņ����T*�1���$�[���Q@�s�G�P_�֒9��ѻ�F��z��>p5ݗd\�"N��i��򇔃c�������K�|�2������I}�����O�:���=	qz���+��Sw�(skh�C܄�P^"�:q��|���aX�61C��VL��k󾦞i6銏�a�س��Ҙ��.\B֢�Z1���h0Dmn��u풇��%��ĮY����1����:�Gx(y_��P/}����:aiIh��a����X�K�w���C��4�\H����!�4nڿ�&����'��H�v�_9!�$��� 燐¡����7��Q@</�Wve�t��4>�+�]G�^�
?�ϫ�+V���q7r�v#c4�<ؗ�!�d��10�r:!љhi�*�1+����A�5�q�����#3 �����M��'h��I(_�F���I�%P�sH��EO~W��D+�?��.֊�m&���z��n�qn�(����@���b��%&^*��[�ז�q�(_�y����Σ�Ã��y�e�E9�9T�Oa(�P-z0�(ب]��3�<z��'��f������`�$0�D.��'[���C�v*���+���J�1��ʳo��O�u�d�ث��!"����=vj:���!hY������,�HG���0%���O? �� ��Zi�4��;�B\@^�[q���1#��a����,|�2�b��?���:��@X���:ک� ?���C�Z���8���H��{\���k=pɎC��xm����P�o�.߶~u�8�D��a� >>�>�PӉ!;����E|�o��ų�P�Y��>�XL㘧j��ꦏ�O���!��,~�_����ǽ���!��n�}L��0�y)�/��~�?̂^_�ֹ��++��W�8�i������`5�����;������[��]Ú�����]��;����7��yS���^���}~�-|1������DS����{}�n�ף�cԸ���^���bڠIQ���lu��[�-pƻ����z��Y��Ee�3���W�,�/��O��=�y�/��^�cS�*?������l:�������}x�}�a���~���_?������u���x13�ȏt��������V�{���������c���d�ח��Kj	h���d�^a���#����v����Mk��Ky�~H6����!/)�g�į��Ǽ�ѯ�S�h��O�쟲�R��_A��"�d����c~�O�¦�lO�^����R�m���A�C0��=[ }�[?K�lTH���C�� �!oL��vT7������<j��-�y4,���E��ӻ��gx��w:_��ϒ)K�Wc�C��70�gɔ���W�p��MR�
Z���ml���?㤖��~r�ؘO��k�l��{�[���N��<������b퐑�m��̖L��s�'e���P�"�iy�*�ܼ�V'�"���rW@6�.�0�r�P*�Ѐ������(��I�b]*��1 ���ҨW]�!�W����쨱�Z�'��_�ѥ�?���v�g��Ϲ&�\
Q���H�}�2Ȝ/�~@y����e�|��[���b7�LL9b^���"ejZ5�(��y�SK�IM���)RY;���,������qps/��&ó(��E�i�I1C����a����b*d?�����۔rw�2tp;����7O�Ƨb*T<Թ�m/���y6�k���G��Q������K�T�p-'�7"�K=��q͒�OG}pשD�ώ���Gy@�
Uz�X�cYc{@��4T���jȸb���Zk�P���;�j�zՓ!�LI([bŢgC��/�&��(]k��t6ڼǡsրP�'�Q�}D�A��M�ʗ:��Ա��O��u�=~7B^(�i�mO�n���&�������R3��.L �X]ȉ���)lBoc���U�Ƃ% :�S��zRS�z|�C�O�����ڃ8 ��M����.�*`{���uW������ᇘ��B����\��	qz���q��?^W=8�Hnm�yNk���EF��,]/���9 �D��thx���1���� �5��a8�����̠Vش�k������(Z�D�����G��&�6����&Tæ�? -kJ�ն�p�!�wѼh��u�d�6v�1L�j7뎛���O6];��f�e�[;Dc:��&�q+��櫿6�jy|�@���b�.o5 \ 
ʘ��X�J�_+��Y�B$N/(zE1{y3ئt�b��^u��Wop�s��q���W�����9N�uR�l�=3�c^N��]۔|���'_�@��U3t{߮�f��P�D�'+���?�:�I%��ԋ$f�X�09����\KӗU<��V@|�7:�Y��5�ӂEk����޾.b�rvB��w�I���`�/j3��1��O�:���@aYs`���I�P�x�ؘ�`��G�6�nD�g��6�"EG�B'3_
R�Qt�(LWF����a.f x����q���G�l2 mS0:�H�4���,ҡp������E@�Q���B}t�<b�ɗ�1��q�> ^��/&�y��/��3a�;ј��Y��~̞;丆<�O6�?h=��,�R�pg��W�y-�LcmLL�#ǂ��lj��C�meoW�oh37�����l�c��6eC[��å�ߏC5p���x0Ϣ�>��$�\E�~,�1W�~]YpR��x>�Yج����v��ga�oV����	�(�g%�& ,E��=�l��4�C�1�����|�MO�Wᐠ+�t�z:s��g�w�3�Ύ�mv�.�u-�`��:��3�\/y,X_�W�y��o�k�9X��E,����h��4��k�G
k��z�:� �2�����i�o%_��j�m_M~���X�YE�ў��i��T���-D̍U��~V��5^?�޸�y�2�q��<�(����zVbA�	��X� �.x.%a����|Ĕ�=�k݁����3�"�������@��
/������t�zk�NAǷ��8���a�N�����BXQ0_��87P<���@������ �V�"����e�R�B��Z���qT�4!�L~�m�TZ�ך�Mt�k�µd�\Z ?���,R��b�+��y����Q����0�0�|mv1�7�r���1����z(n_&%��臡\* ���4������t1�j.�C�P���y�G����\��s�����X���Pl��$@���oN@�=�E`��$��o?���ӂ��8�3�]*����"�~�q|W���W�������]W�wՀ��8�{��r�y�8J5|�G���4��kŢ</�w�\j�1._����=���@̬��@��I br
L������B�\�}�k��Qd�n��b`ʳ�����k{]J�ݴ��X\G���k搿�]* ���j�i`�u�O�e��F���@����w�m�����1ka��-�=��Z����y�?����O\��"zn_�,���ǻ�A5|UN\����!WL9�����4(��1]	��s1�b��)�D3�0@���j��`�}L:����ѩ#Ӝ���aPԻv�(���v�R�D�X*�@ə$��_��CƗ��^S����M@yzw�v1:���Y$M��c�b�w�e�퇼��9ۋ��rn�����Y?=\�!� x*__ �G��-9��{����U����X��>X��8%��K�`�Ë�?���/K���]��<Z#��i<�R���U��������ņ��2�o��E��Т�>��jyx.����f������o�/�d�]#|��������G��3�
��}�����H�c��&?8�6���ŏ������~�m���K#��|��m??[�G�U	x�Cý߬��L���>������ٿ3��:��5�������@.�_�h}�5�����G�ͮ���v6���������N���'���-.�I�O��[���%
���/�k�!Y�[j��w��2�[����Cބ��~<�m���C�r6��t��9�Y�̯��?���t�%�?��k;�S�g�qY��VV��w��ӡg�|��_$k���ϟ<+����C~��
��k��y/���Ol������?d��>i��q�)����lY�=g�
�����������VCc�s[��7��EjF�7�v�?k��~<��]����=���3�Hp���?-�����%���w���S=�:���ۡwv������D��P��d��X��/*f�]����K-�J%��\�a�H��q�j�s-�T�+b(�{���I��;h���V�FA�6�X�"K- �l����vW��w^M��^^@y ��y�a�+���]+��pcԀh ���2H��\�N(�&�$�0 �jȭ'۴e��Qt��.�Bz��U�KV�ݹ-Gռ��� ~6 ��k`c�*�>�����"�: �����T�g�aq�yѿ` ���)�K�ױ�7\ܲ��ć����Y!}�)tC��j�u�㨦 ~P���B�Y���������P�����a��r#���3���cVY}�a.=��_2yX1���/�o�sŐ�����]+�ӱ\Fm3x!���Ee���6��Eg��9����:e	aYC&�|�j#S�6���E����b�*V@�����T;����w,�QGO�o{ ��]����T6� �-W��_�V�.+���{s8�z^8�W�1���'d��y���Hﮁ�u-,j�{�u�׮t���p�cDCx��C׍�K<�	�kE���{�=ԣU�O�������Y��=�`ʍ�nnr�\+P��&���N�����G!<��ݪ*�8�!�#���"D�Iy�3�f������u5)�s�8��N	�J�����L��y.F���[)���C*��E���6P��Ǵf���P��i�&���x)�@L&$�6I���6�ͮ9����^�|~Ћ��K��0Y��@%}&D�\���EBO[���_�v0���U����n{��d>��<����Z8��Ƿ�B��4�w��밋�yrMC��ky��v?�Z%��k7o�2Aꆗ�g���������塼�� �0�w�彲���v@��+b�X�#�7�W����= �W�]+�Ɗ�7� bP@Q�Y�t��WX����ܥ��/����,����c=1H,��l��ﯭ�G�iT|z4���f���ܤ�J�UV^�)G����g��T��^�h&������]K����->��ڛ��*����p���Rq����S��Ї��딖������+�}����e�"E� �]}5������5��@�\�>�!�oB�Fe��U1UN���L1�"*�iT���IͨD���E�h8Ĥ��^(�=���/�<P���8�l>W�򳏱)_j�y���y��G�n��õ�H�`�n(�(�c0q�.�FH�G��F�c@�˂�hח<�Y���jL�>w����ܨ�'�;<�'�S��"�';,�V,$`�P��{�c� 6z�)������L����xU��YH�����-����(~~j~^�P����E@�|#,9=:��z�����U��_e��_�,4�Y��-xdH�we�s����+����4\u6����\(ϙfc�ȣ�����������iO~�IU�{���S�+��Q�w�w�� ����+�G6ϴ ���LK�s0q��Jl@<��"�?5���~�6����D7$����=(���̜�$�C(o�ͥ�<S�k��j@�,�y��y`�b���6U��r�}����q��'�C��`�<��<������%��\@Ώ����Ķn��ԇ�����l�����
��*����;�!\��ejƪD>�J}�BH��\����F�:��r�1�R�j�S�Y��/ l:V0k��
#�����r�> ��.)%5��DÜ����8z/�!���LLDi�����ᨉ���`!��f�]�F�x-���۾�Ob�S�F��Y�%et�<��z4�G~�:ۏs�\��Ӽ�?�߻��t�J�~��b�����<: "�L��Ĕ��e����+��]tvĊWe[5d����W캮w��Rۓ��nl=m���U.�A�ڭ�tn�xc8��>��n�������I�]Q�C�L�t��l�?��n4���x�yA��J���ȫ����:���|��=U�Ol������zh����,�CW6�޾�o/z�X���\@<��n/z�Kh���pڋ2O@�~S��n�����ӛX�܇-�+�TIO8T�l�9�<l��t��(>���J�|� �q�P������lH���Xw拨8��:�CWܤ�ѣ�oHnz7G�kr�t(��ӺbqV��ڌ��8��;CA����"���Ar��W;p�9�ݯX<��kK��JD�ly��̑����(jG^G@�,H{q��rʉU*�JXL�c������!?�5=j� k��X��,�|�wB��2`-�����~b�<=O����]�s��s�ֈy�>�u��!6��#9���>�)������C��}d�C�5P�����]�G6��|���i2{�K��j�wU���s͵+ծ��tW���I�L�������oz�m+�o���7u^��V����y�R��������{����;����mA_\߲�����x�?��>�O��G:������|��Aߐ�ߜ�+��CN��~����ϑ��L�W�����2Q�|����kj�I�?\Ť�������5���,5����S�y,Q����o�����=�_{�-�_�z�����o����h>��c:���%��#��9<��]��.�)G[�"��%�W쑐��'vo=#Y��I	���g:&��$n5���)��
��}�����H�O��?��g�[�[}d�v���,_�O3#/I�l�����g���s������M����1���,��d,���,v�
g��pr�s������s�zrX�G�����a�l3��-��D>�
��M)>��b�w��!-=�O��?�-���u�wm�C��)�
OAj�j{~���zO�O�Z��Ȧҟ�a���E1����dM�+띝qz�|s��"�1%��y|��(��.�u���^�"�B��T-�+c�P����ei��'��굢+��oQ�x���ph8�^}�Ԇkf,e����tl�bN���2:3Ԑc��b.��z��-J�"�}L�*�2HB+�<�2�Ί���Ɩ���X}�^�Bi�����/�x\4�.�p�vCF�$#��H���P�QΣ��ӛ�� ���r�>���s��Q
6�mA. Z�.�Q"*@�m���&xs��];�Ǉ-�z{w!�����X�|���jac�*�9J�+B��G}9� �R����+ �����ZM�nLb&�ێ�Ga��T��8�A1 ��mr���O�P/����9
�B@���}�i��s+o�֮~(����_�ӏ���z��bȬ� {j��0��v?a��e�]
��?�(6hoM[1y��K��b�ܸ��|�yH}?v
GS�����!R�f�-��-�ŧ��SH�>�"��=dF\��|���i��㪽����p�́��39��*:��
�u-\We���W[��v=���u5qʭ�]I{����?D�=-B�N,U�l�̃��u$�B�;PT����c���'"m�? ��S��I:^�8���L��f�t��Mϧf�]�p.H�mM���X�u��j�6	�� ������3����0�V`!T|P.���G@y��	F~�!�,h�b=a�7 �܉�� B��!���^Qp�
+�@�A�ċ��"��굱�%�v'H13!w����a��: "�u������4#��}��Ѿ�{�x��ģ����/�$�%e���p�y�I��yE�O��ZD�$�l7�I�a�3��
�%�a�����!�z+�?���Sx8��h�b���=�Z�����(�{X�g��{�d}T�=��QX�\(��`�x�x��z@hP��X���υP�><U�GG,F9=���SXz�L����Ѽ�F�7.@74_}�%y�|N�P�5�^���Awx���|]E�PB=���𪀈����c<u'�9�
�R�_�z�wQ����9���71�c3��oh�p��R�5�<�cF���>�f]����Gb�A+�<���)h����Q��0y��,+��
;�L�y�9S^欰�g5����yct��
��78x���>{����fexu�(/ko�M��Nz��ة^�f~8ב9X�A�],��%O�V7�8_Ĥ���I�e��ui��;���{@���s��c)�]P�Eq�&��NG���:6���ڔ���}<A�u(#�
�hp���&(���zؠ��5ʸ�#T|�]=#��KK�����4q�T)䯖����P�{P�uS�QR�PX3�k
��D�
��R�XMuic�7>��Y]�d���,b�������f�a�� �����Do�Q�5n$���$�,�֬4���y@y�=�jIj��C�h��b{m����U�et�'��Zd�1%�{�|]�H�A��$io��7!9��Cm. �ɡE�G��xB`�ط�{�Yvg�\���<�̍��! . $u�����,�b���]ՖU�62m3�]��h]����k�s-����ÕR����\��-�-kT�B��҉��W�	�.�W�m�������&_��rϴսo�0w�#k��7x<��PΨ���\�6G1�\}&�Kb.�P�����#UfI�1I}�P����ٞlv��ƞ6�����Tř�Q{��|c�9��=�\ڋ����2��q���U�:�ޛUS̆�Ko�,�(��'���дCy̿�zRP=Oɍ��~5��,;*;���1��P~:�S�N��3��:e"A,=X���|�Nů9�0��*�E��DEc(z��/_@DŶ���y�i��B�֔F6���A�Bw��c�%���wh�F'�P'a( ZΠ�rե����3��9*�τ�v&[b�����2@|��V �G��7��l>_ѣ
Gf@�����8�\�ܛ�$N�{<����+?���9Sۇ����UxW�=���-f�`�5�x�w���}6쏿�Ze|�`/[���������CTX~��ox���ߘ�x\���ifmL���}*j�f�`�2����%?|bh_]�G�7�P�=��;"���|�t�5���s 㒦?�o����ȖX٣l�_���������u������@ޚ�����L���N��������?^ǧ����w�O������}I�׳lo���Bvj������z��$/'���yv���w>�"Y����6�m{�շ�C��ԣ /���$�vf9�g��|�^@j�9�"���VP/���NǓe`�����3�̉�=�?�dA��Y�6{��O��O�3|�+o���ם��:_��+�K�n�,P\5�j��V�$���E���O�m��1�~s�^	\��}��q�����9��VwH�>=��@��Nm�!3���_SL�2r���p�
z����I��3���z v�\[��*�6*�R��Q�_� �2FϬi)���f��{�o����s\<�<�'E'��	�b�w����������v�Tކ��%� �3o���oe]�V�[b�� �$C>�B3B�匞��p����MRon��7kr�ߨ�|���,�e!V��ߵ�h��B]�|�{�ea�l��^w@&�"ɺP~�-�rL�qN>WX�����XۡWS����{��HبT����1�'ݯ�����2�_L s��r����$jGW!c�
�5 d.��û�2!ӢBU��̥��u�B��Q��_'M4S?W�����p�
��L
�7�$?�9rg��<����:7J���o@�.�c�G��V��2��\���{39��[u���Ϻ�Ý���z`���Ш�j�tc:Q�M�B'���,.C5�|�,'yH�Z.~8H�{p׌6�KS���&}��~�MӂV�,Q�m1�BFUa�����l���0(OW�O�j�W[��5����w5Fb������d���P!E`�h�x���A��A��L�qI�yn&����6����J4�+�	e#�6�TS� ����p�o��Lݛj�6��'T��P�M39�!�n��凳���<��Հ�^�G����y��סQc|y���v0X%�a�q����<׎/C9\�19
Q�����0����%��k� ��z. 2z��b����ﭠ�kđ��ڮA7��1����w����\�(N�3�+�CGg�XH����A5��?��鑓��>�-�s�ƽ�
e2�y���D��XI����]�����Ă�� ��5��7$�����p��#�k�Ym\�����7��}S}�:�|C��_jl>�!���!�#�a<���t���w=�hM|2.�ڎ����:F�E0
lܡ�����Q�X@!w���%�o4��bZ�^���3$�p���j�2h]�B�<>>�?;��)ݼ�o�N;3�#��Bl5�M�(ĭ���L9\�M�j�X�̎��$7=0C���:G�	���|]sq�U�x�v̐�ZDk��GT$�ō�����Ɗ�
�8�$Z��3䧰�č��&>"�#&�B���q�h�^.k���sBT��O5Frr�
2�YX��xoz$�h@��BYU�����!����P��`��ʜq?����F�k|h������7Չ�۵�S��G$�::\}_v�޳c�7�QxH�n�"�餃Az��3b[�򙳘��9�'�~A�$� �B���Is�*�<ą�溺�@�L�]Ԛ��S�`L|��N��DEn�b�E������J�U1��o$c��� Pn��a�j�iYQX7>C1*�B)k��U謮rO1�EU���
3�Uv~����4}U�9b��j��dr������Yw�er�j�~W�ci]�u���	�	�j�6���jp�Wc��B�Y�.�p� J�2��K�n�s�@�?D�{#��v�ODGKx�43q���A�j׍G��& d��`�E�a�C�����-'�����c�.�j.�yfpb:Fb1��:,bס^��=�HF�|p1Bt�0{�۷��� 6>*��X&_�|3�����C}�.T��N_�9殅\���!uaͧ��8ۍ
q�9wkQ�'��m���}̀��j�:{0�P��1��ݷ�G�w��u�&���zl(ExS��d�&+rT�ơNv��L�]G;MћD��u-���]�
���_\i���7[�7��sMћ���Bm�T?�h=p.��ч8kom����[j�Rsm�w帵'GY=<��<���`Nt�B��
��W��Q�B�v��<�T�b�Y1j�U�D�+��H�*��ט�F�]�Q�r��:S�c��hv��=�����;�Q����BmI�~i0��Yh�O��Lxe�d?�B���>�rp@���4�,?d8g�{6^FW��&Ϗ/��|��#ʌ��\�����̱�Ʒ�����s�3<�FJO��ڿg����Z���~�bSMݳԘ=K�߳���r��?~B�+/��Ϸ���C�V_��3����0C��0������n��������
��湴��mSe{U?�z����
��}�����������~*�я�e�/��<�Q}V�`�O0a�>F���Q����Q�?��s�K�_?���?2�+{��P�O`�ue���g��	J|����w꣄|�m??�KD��Z�Ov�k����������&��^�����']̹e/���Y����C��j@Ֆ��n�FB�Ɲ�h����3[�	d���Nνk�U�?��;/�!���Y��Y��d�Yy	/ɒ��5�NR��L�YY<8N����5�Fi�s�l��N<~9|%#%K��;������k�vn���e)�n�
?�Q?�`δ�D;�r�������ŃGS����� �Y^|���=��/�u>����W��eD�Qd�C� 6rY�{��UH�����ʢbBWQU� ��B�s;������h�]�c�O�[3��%Kl�ï��q��:���q퉅���g+3��:{^7���2����T�unh`MJ�IrE�l����!7옣`B4���m�`��ъ����i�R6;�!7�T�<`C�(�A5x0y�������Fut|�,��`u��������Bc��Q8i�b|Y������=�9h���GY��v㇈K�������oj[��N���PSwg�!z�2w�F{u2)j��Y�+W�S���ڑ��n|�P!6�ojG�X���F+7pӮ�H�j6RL�ФMf
��'e�X��-l��R���P��e��f�Poy��<����">.uC�����Z]D��DH�~v=��g�	���ny&{ 66����B��/����J1ȭ�YZ@h�
��]�1N�FX�G!��8j�6�h��u~�����c���U�Qtn�P9�����k���Ȟ6�V]�[��g�Mf�m��|����!|�v	d	ZЭB�f�{���V
q@|
��=i�Na;���yЉ�=O�@�돊��L����+��0����*z-�g*3�^W^]æ�"iLz��QuA��Z�u&AvŔ��a���bf؅�p���.��J�8��O@��-�?��xT�����+4C�̦��B��0�	(�O�e�[��*?�]�BߨRo0�$��	ݽK����5DFD�f�.�K�01���C��B�\F�\itV�4G1��PD��B��r?1*U�X��1-�N�k��� �iM�C�Z��Nü���Iqc<*xLZ�s��4�+�ǔ�	�iL,љB5�`�ɟ�bИ(\���!x�5:��"ct,�c��5n�C�`��D�t���ʊW{�O·Oa>�Χ#�x�CMg���Bg5��W����sU�g��> ������X-���evW�hs�<^s>}Gy!�-`SN����L��B~ҡd���(�+�!�A8'"�9�L��]G#!q���k@�(�{.�ѿp��(��K��ܦ�m���>G� �»�  h�1@��]��Ux��9y<TҘ
��U�8����L��#�K��ai<�*����Q=M�1ݠ[��F)SY��4��py37^
E
rÀ�(4���ǫ��O�cx���T�A4Ί13�ޝ�5�U���|�ӿ8��\���Dp��Ù|�k�41M�P���3��<�\%1�&Hk7<����H(���m� �X!t�hF/�<�O�=�U�!�@����9y ���0P\3	��Zi��r�'T��ի�j�ɕ��g���Km|
�x��2.��ܛT��!o�l�������4�=ȧ��_5
�?�/uȹ8�d���+�=M!�T~.��w�^�/bb���ܓ����jOX���dd��¼�Ffr��p��7�.{ǵ1_�fD@ė���B�qW�s��B|����	��_�yP�gr��R�䙧04�l���
[��R��jnP=�[���q�4ȧ#=�ӛ�y:٧/�:y�G��k�8��(φ�@?y��D�Z]�A~^Ά�0Ai�<4�Y$P2:�ę�َjwpϯc��m�J�9�\u�4C�P�5Vg��(�q	�bT��̳�c�e@��H��t��-�����:뇖�W�ϯG�P���W!����F}K�_���?��o�����?bwF�~��-}��k�t&�(�݉4�V=��f^�q}���=D��E�?���x}���y�m�A����g.9�e��܇���->��ב����cs�6�������lp2���_���H{22~��?de�u}S���t��y�?d���R�ȉ�ͯNNuiO��仈	r&x���7��:g��E����+��e�d����>J���~HNQ;�'����� Sһ���Ǽ_Ë�'6_��;����{_#?�52�}�|�kg��:Yz��0o=�G��E�5r��O���#��y^a�?��k>5��.FB�X �\��G����}�^�U��pcV�h��VnC�*;0��,sU�R�~�PP��0.�:�ņЅ�=?�x�k�d �mo�x���b�ɻ�w��W?�����b�-eN��j/19_�z�>M1��,j�Ű�rS�P>l6eʆ�T6l������<�ͤ3��}�J�=�L/��Zfv�k( �b�M���o;��T��S}0 �I*�wzѶ�AP�T�N(@8k�B����e"d��B�a��*ǵB���Y@I\�U�:{w��#1�,d�")�{T?S�t���0��0ƃ�V'�Ѕ`�Z�!?|�"���EU��{u���7��� �Q� ����]�CVU�z0h���q9�0�Q��D��"[��j�v5�@�Rci@��îI{��I"!���9���po������_ ���t�XM�/���
��[g�rLjDe �5���e��7'���+���p�|�I��`�[��U�O�z�gh��6�j��6��orl��۞C��"�dz�!ۢ~���Ɯ��2�ED�h�6�fS��?�Ҿ1|j�	�H�?<&v�Flȱ79�g�|3�2 ��uQ��&�������~o�/u#5�E����i�  t�Ԓ.��ld�p�#��tH(�P��+m����m��n~qcN�52�6z��* �P�αw�]���u���m�ѣ��Z��i@y^x�ޜ�&7v��1w}���S&��0�O)�G�.�O"��r]˯vѹ��a����%
�Zh�o�G-^�2�e?�����oLݯ��H�rN��.���W@ҽ�:F�Y�f_gVm�k2۷"�FE�f�����1�{ld퍆w��8s��P��g"���/m���f���p�^n�E�0�_��GO2���!�d���P�7�������2�i�C?���}�yOu��7�h@�l�C��2�e�&��D���L�������H��Uv�q�
fi�Ęs9(�d☒Aig64���������
�-Cxܨ= �g�aހ�"���ET����8��睕��k*��]�Y	f�T{΅�j@���y�W��:�� �ƀ?5��h��, �j�gt6���$�`Z�g�1�wn�!l����WN�QTEb�E��f�@1���0-e�q6AKѷ�I͜��BE1���B���M��sN/�YG��i,R�w�g�s!�Ȩ�宀!�k���q����<����!s�{���f޳1��p�&��n�2�r=����+j��׃�k�,
� mbUt��(*�J�g���H��@�%���Ѐ��":@�����F�%�Gy��N�2�=ֺ�=�n䁒�y�Ng8Yr���*0��K���qԁ�? h.�"W�>��|8�P�	9z@�����c�F^����,�n
F����ƀh���|5����m�TrH_�&^�A�]�^��
;�4����HA(��_MC>}��+zh8�1+ȗZ1u	���LNwe�ߕq(�,����v�n��d��nЪ�������ڝ_6b�N4 �n�*B�07AX���� �6��q��1(,�i��$��/�d�O5���4a�a����i��
��k@�@�xov}�&m`o�	� �-�# X�%R@����Щ�A�AsP6�����й��b�r��Z������y��G߰��T$缠�9����X�����x_!�\+�|������O�,b!�1>t�)�6r�q�1�4�S8����4꘍s,��nC���D4�kP:��3�'b�@l�`��D/�,���Zj8�(�X���;F�A֙��b6t��7�:?	����-C1K�(��Vu�!q��������8�(�=��O2¯9}��B\K|��� E�9�R���t�//!������V�>�_w�b�x���7��|�����;S޽�O����:u���T�[=���w=�IP�Y�����L��i��7t����Ы���*}d#�C��V䓖`JC_�����m�Z	_�r�W�����>ƻ\{�!��>9o��+9o��7r�7/��K�G�W	�	Qxǅ_@~��?�ɯc�#����P�a ��^k�Ԏ���
�z2���h�~���	�O���'����"�����y@�N~����9T����A�0^���������!Y�0��b���������:�|ͫdC�5�t������j�=ә��ʙ��;=?��2!�v`@P��J-n��B�SѪ����Q(N�KYx՗��E�s)����B��K]؞��_���8�8opxK�}��F�w<�?4�Po��k9��5B��g��,8�ϊ}��<��	y��qU��V�b,�$�LK�$e6�eaz\��{�ų_��ͮ��'�L�����C^[��BJ9X�FϏ��l�����i@��	���$�і�!E��k�ȃ/R��((خ�U�{%o0>�����ph������P*T<���j���cr!�6uͧzmv�)U�dk�دk���������:bՐ	o��>0��]��4��u�WAm�؀T,B��f�:.��q-�V�׺)�\�*��'�@�t��VC���eI��%��I�!�1������7���+�a��B�����c� mCͦ)m+�����iufV��2:BBK�`����Fv�'���U@y���rs=�h0�5`o�\-)�e�6�(ݞ3yBH�P�00 �'OW.k=��駮�����'a�؎�)B����h��(h�b�[�6! ���Ų��0FAAnǅ�Y@����y�ը1F��l*t�Rzy��K�h�'Vץ�;]���+�[��A���m7����O/�7��1��њ��i����W�Vw�#_�\��t��p��m���GA$0��]�<G)�0a��{B0�*��tǇ��'��A$��{=D�%x�M��B�R7�	}Cw������A;��+|��!>(�<*�t�sQT��Kw|)����l�gA�V"?D(�9�Aߍ:=���.�zVd���a�Ѝ{r�n�o��ʸ=*����g\Eq�Ai��e4�}�!{��g�yg:<:�w�%ҵ�G.�2�z2aя��^��H�1�2�H`BZr���!�R��0)���R/�lrn�\?~�����r1�����r?q�|zM0c��hÜ��{<,�����DP#����BV��iy�4���|��ݙ�\���,��g9yT�p����+^@p0s��B�Į� ������Z��O�l,<��� (��c�|E��3������b����?�SY�$�oN���Ď}*��o������Q��N��ϗ�,��c�%���-w0s����K��S�6�0>� ��5?�����p��Du<8�Jz'���ٱ�gn�n e�fkWepÜ�ET�:V+����հ}Y*�5^�(z���Q�}��Bg�Y���]joV��bޙO?p�2����K���n)dh ؟�v�����n���?��  �e�2��~�x�S�(O���җ:�ˠ�#��l �ױ�7^���&��B�\ǿx��9Evj@��<�"��PtYn+�`�L�}t������]9���+� �x\��s�l{ֵ7� �>���*t�A�.h�w�U��m\�=��'wi[����+^���;�h@r�Y"���qwV���ݨ��|������p�������{aH�ojN��D�b�:'(���yz��7��}��t��G/�i{|������p��I՛��&.fZo���r���4肙a@8�W��+t�6��Ӆ�_��\�7��F�:���}{�������1�z� �w��"&�ˀ��LTHіxSb�d�y&��'&�P���<+�q*�ӂ��I!g�Z�N�6�bÌ8�������� 1���>S�r�8�;��7t����#��[���K�-�ׇ��k�Z�4��c��`�<_�����������m��������P��8��{��ߖ���ո7�K�?�{�oU�K{��ƣs�(:�w��О}G�����5�y���A�G��<rY���~��ϑ�?t#��7=��c�ow���]~��;v�猥�� �M"��f�D����?��_g��������79���l�^0���E���L��x�k�CN�����_$�����kn���k���yuW������1��mg;��2:H6x�5�W�P�{~�"v_�
�7a�%��Cn�)!=��b̑�w:���]�虀?g�oϝe�����3��|��Ϳ״?�7��μ_��i~�切�:���t�g`���8{�7xp�*�M�k���Ce�Ar����*�Y�e��e�gFmek�����W*0��-x��?p�[��(<�'P1���-���5v&JGe���һR�X�?z^��A,sĭƐ�w�ʠ����z_n�	�G8q�m��V��ү�<��A4�f5:s��}xC�rP��<Y�)����2��(�~:_��2�r8��r���ھX�σ��_�>�02VgLG �>Z�?XG�c��`rP����l����? (�f�_j�<x���ȑ��FhK5��Z��7/y#�����hK��t�����g��k�5+��V�,���&�fJ����(�x�U�O�����8�A��j�N��yOC��ٖ��7�F)$�*yՉ�1����y�%�P��ƅ�*� 㓡S��J���[��fD��~#A���z�l_����Zg���zP�q�"�7�?��7��v�T��J�1/lR�Z�v�m��P�Չ�
�UX+����O��^í�mߚ�֑^4���}�����U�M�0�^t�fm�<h�T\)��pC�o�I�MBl�n�M�����Rp�ҋ�_\�OaSl����Ѷ���CüI��m�aR(�v�ٻ.=�T��C�-D����<��[��+3�^1�� ������scm��?\p��w��
R��(��ѳ�� �M����0C�j{��x�1� Q������	c��ohl��!�`R��6����~4�}��0��U�<�5���MnA��S�~�2a�{�Lf�� 6��?�O��>��\�6�� LwcQ��k"{�x3���g��x�G
f�C�x<Z�#[�a��V8�^�G8m�<�Q�ލ�JdTVұ؂R]u�w/-�<��n狨���g�W���)��O����p�3:�#!"�0�$�dv����!ߘ����� �}��7����\���b����|8�P.nd|�����&Bl�#o� �r���= c`��}F�P��G��G���h@�y�f��"��H�Ec�rp�� �c�)WF���Q�k@\jÆ�z�st�i^ʔ�r�����m�_ggGdv�}��*:�s�1{S����q��"�tfu]�9��=�^�!n�J��.�|SaR@y3c�-���d?g.̓/�b?�����Ob��0��0��p�^�W�D�!�<�mc�J{��ЩHU�Y����@-���
K�A������p�a����C3��y���W�:W!�a���0*\!D��Bg�
��UKޏ^���l���d��=6%!�jR��S�Q~� 7��qT���E�6s&�Uru,��N�}�|ұ��||k�����z�
J�|n�lDPX�`!9�J���mbSY\�r��5����o{C��f�h#�u\=C��yh&���ȕ%`�t�Y���M03T��D@y�y?��?��oY̬�u�D�R�D���&h�+�ͻ���7���6�R��)>����+�]Y�q�6�/�h����-�A��̳{����ٵ���Ia����l9n�]�~L��A��Vޠ�G�}g@�GM��2�bѹ�C���T`A��2�M�< >��H���V>�AY��P��̅8��$�W��r��	�p����2�:yYs�]�A {�Iʋ��.<���WLW�PPxS��J�X�����M"�\H�/��zpJv*���tz7N���=C�����1�zT����BVu%!�H�t�C�q�t6Ib���1��r�Hs�I��Ԙ#/- �q������7�����L�����#�Z=�۱L��kfx6ōrS^�_܄�\-	� �E�!2V�����1�R	��a��*��a�U��)���.�����y�J�w���D6��?T"������.�(#����Z��y\�9���U���:��olC��9�?�"z�C��g�/���un��g}�]s�X|���/�[~����L��%�G�w���k���M�x%�ݽ�JO��X �q�����ww�')	�}��d"�[{e"YR�,�#��!����L��_��׷��C�$����sd�����~�ߘ�C2�?F�$qh#��R`HOH�S$ -;����c�w�'9+��G��s��r��
�����>8��2�[o
��op�,_X#t���9�1;?����'�qv�R�]�_�	HG8�.�H���[�>Y,uj���T�sԒ쟀�������C2�c�����";�޼���L)��_=_�*��7q;�0�\��+�|���n�G���.�9��������8ܖ��|"@~VPe����� ��=��&�L����;����Y�e���ϲV�@��F�3���O@�4��oĔ�P��1��~cZ����7��빖��h���ulh��M�r�Ɂ�3�ńI��ݢ[�F���xu!(>p���³�/��c�s�8���
) �d�W�����#���Q�\>��mZ��
݈�~��_�U��j���:̀0m��+̂�E��UC�� ��.��cj* 첛����Ɵ7 �:��k�c>;)�Ъ�~nL�a��-.s�Dހ�"��|�պ���}6�[�E_ɹh���ɳא_F��}�W.����E�\���I���;��qo���X��6 �3��Cv6c2�Pܶ���\*~gm>p�|*N�L1��=�����]"wnL�*1�����ffqtx�˷�m�VJʛ��L�0o�v��t}���P������1�����-���^�Ѹ�up�o�X�`���O�:�W&"7�W=�����7���}{��=>6�3]�,���~ӂ9�ya�	Į��Q\}� B�棉���I	,&0���T�O��������h_���}ЛЧ.��F�r���[��&\)������]ux?��b�Fd�Q�s�(�N���1]��6�T����~<��#�b!͹
:�kȟ]۝��2��d��Qh�7��s�I24�2G��74��v/�*S��>���0�lt䏣���z�����02N��`й_�~������7:N?)��ɸ=���~�ߏ��_4�#�RVc�<��^�>^��A��$��4��Z�f��Ý��������u�SʤcF�=���`%<N7s{����U
 ��3o·�㴳�;��V8��Y�R���kȏ6נS<��lM9��K��_���\#.�'�j�D�Su����� d���:z�ّe^�?�:s�ڝ�x�y�r�a�ˢ�U�Ԇ^W���ϧ_���\��'�m����������Gi>�A<�ٍ�\{�;�}p�U ��G_�G��[<������k�k�H/r�����v��x.����3'�
����0�u;V��{�4���S�5cĄ�`��gCk"�_��L��dg>z�<�ư-+��D@�������y-��&�蒻�um# >���\�Ȅ�֥Q�%w�0�V{���6���&~0$��4C��o( ��_�=>�Js��*�����Wm��� �ׅ;���k�I�Mc�Fg�m�5�鍩�n�կ�C��6_�7���{�ow�QU^,D�m������%@�&�tOl��1{B���|��x�kC�{�r^�|�up�_H��1�aV������Xx�:�|o�q3��jL.�;��a�?�<�]�6tr2=������8;��!��:3d��#��aG�<'`�Pt���By8�^;��S�v/̬�y����B>�54�(&H�5̩��YD��t�ף ��BUۂ+N��qZ7�9 �}c�{:������թ�땒!��4ڶ���������W���L�D�u&9Pg��:�t���YLO\|f�o�O�i�@�\{�L�Z#P����T���9z�?E��ze�ؔ)������~�C�`�X�]ޚ������V_���M�/��k�/#��/k���0�iy���k��2w�����yYM6��9�徥?�5�Xֿ�͏��k?��Y���_��o���a����=���'�Q�k��C��zt���F�������8������N�ee�p9�̟@��ԫ�.�삿���ǖ�d��ǧ���Ͽ��o�����e�m{�	?�s���<��|�d��Q�y�ή�w�1!-S��xVF�����Ε��|G����L�y�L>�'��;��u��ٴ������\�g�L��o��ϙ>���u�ɶ�!�K,.�2̨�+�HP�(8>zx�����ac�9�A\�d ���,�4j"���0F1�A��,Jx�w*e`hé4a��� >�v�� o�(a+Rq§2�(�DⲐ��V�	���Ք�GP^�_�+F�VxF�;�G���i���Sk�X��]׆Go��
�S��&�����~p8~K���u�T7٫���5�,Q�x���8��J��:1٪78CJ���ui�}��3T��5�/�u������3�0��g�\�$T}��S�U���L����AbR���EM@��>�T_#�L�{�\�A���Ik�j�g��(���r#���P�����j���f�p�j�E4��k��b� a�n��Cn�]��
3-q`�L�l��6�\6&MR��P���K��s�����@R%q4�`��N}�����r��D�鹏��M٘̖��o�av=�c)�Q:�VYi�d�h�\}�{�	�~
��]�t��R3��N�%������Y���Ǆ/;�V�˒.������'���
]r����z�ҭ*D��\����m��ـd=R��	��MY��狸��_6T��c��0�]�!\?��C�(̬F��0*����J�0/& ��e5��e��oϭ0��X�@��qx!.���6:�&C���{��&�~�C��1�X���l0��V8f�9�c���n� �������R�XD��Ÿc�s΅��X��������@8$�6*�3��/�7H!~�/#�a\5�k�7�c�,$ҹMLm㦊�Y4��~7�J����l�����j�Z(�DS��> ��Vhc�Ь�_g�!r�8�\��l>�v2U"zBL�;��i����c͝�e�h5m�9��I�ۜP^�Eyʳ�R��:�T��t����|]�lɹЀ�ea��_�&P{n�7����	���AH#ѭ�z<DVL�z� �_˖�z�V�,zm|OU��iT�3t�Ȫ���ppy!�i	(�ᜋ��u���3�q���,�ʤ��١��#lL�))k��O� ���X��K���ȹf�T�+
�J���Z�'�f��웬}������+�pxX���8=^lѡ�}p����݃p�C@��{��T��ץ�pK����.t�� �f��ޅ��m��{͗Z��=V�p+��X��n0�">=�W�igL���z�B$ '�Lθ��R{��t�����7؅�X��|�҅�97�v�5p!}b�F.���J�}� 1 ��bδs������l�&K�$&
m7�*{k|��^� \?F�X��U�>,��ac�<���ݻ��õ�	��5��������>���e����) ����Gxk��0
HN��0&m�K����"����� ��-�mU�Q?����B�k4�A��l�\wT bn=d<-�'�TW�o��*��!7�/^�K�Hp��W����A-_�n�%7u�Ad��ގ	L�Y�*-'������UՋ�y����_�����N?l����V9��ʃ-�s�O��X|z��׺��*c��ڈ6y~��{��>��������u�\�����ѯ��E��7�oL[8_z��?���,���3o������$����1E}}^�zc�^�b̮9g{^�������wG�c���}H�o�����2���u������U���d�\�&�1��M+'s�j���2x<�̬lE��lZ�����R��@�W�Q[� �����M��!���d͏2��.��]������7f~�cf>��:�������n�ڗf�����X��cx�}��V�iS���{���A�W���f!���~f�]�X�r�/QѕgX%Fl?��U�ъ�u5���H	���b#J��	���ٽ���Zi��d�e�2q%���x�I=D�S�~�����(@˛��ILg@z��V申�R�L�K�DJ^��]kH8����'d��I_+�4ײ���B�w( ���
2�=�+y җ��$��kՙ�1�.j|}�wb�T���
T��90\��R���j�Q��yb]�#l����uk���Kfc�6|Ǯ�M��
a�^NQ���v�=U3�Kc��~`���:ؖ��������:���'�uN�Br��� �kC�\�yԛ����7�)5F�� ��v�1ȴzh���_=Tkt0�7��l�sA �$L�����-"�MV���叵)C@{��,ǀ���T��1+��3���mG��R�PfIV$+Đ��f\�r(�9��uk�G^�]~�:w�B9S���,�ے��ȡ~i��	��Q��0��|ڡ��AqMA�aBBJ�ӕ��|�?>$��g塩D��ӓ�����߯�'C�]�n�ê�a�Z�+����mw���jNb�۵��Uq���JW��;ax1e�	4�;_}\���Uz�8�v29c$��B�����unLr��/�-C�gv+ؗU�Q������2��?���V��Q�t$C3��1́�K�|��4* ��K�n�i?��)g<pE�C�-�_yV�������g%�S�d�U�bf?��>�Z)V]�K�ՠ1VQ�!�	���'�a��be�;�њ<��Q�B��ౚP��/{$soW�!��a�s�"�8 l,U����ȵ������:YH](_ל�EΙ;���ð@~��:nbPy��3Dgu�M����]���b*���$��A�:u�ڇX�o�y�}2T0#,�s2H�b�gǲ���8+�ٞ<
�N-�gî{6\��u���<=��S&�l(8b�)���:?n?�gߵ�h�6��Q��VG���fD@������txN&�N�`=���{.���
���kv�Q3�u���6��^ǭi�CC���֣��3��{a.503���qA´�����/����ifV�gr������K���`�V4��c��u� ���ų�ՈUZM��\�k��Y��7���V�q�;/�вL�]�V@y��ё746��C2���N��\pO�b��(�L��<�`֚Zu⦻��Z�t��a�f�k햗�kw��a3�zSac�@!�VN@��������Q�\�i!qf��K��Y�6�X���h��~W�r�2�(olܵb~�����tw:���,vR�v��9��%�>±�P�}��v= ��x0����ųc��A%N����~cl�ْ���m?р`oF+�T���������ڇ}���=��P����?�sʀ���kL���{�~�¶�)���Vʩl*�=�|]M.ec�|�K8
K���8=�wG��qU~��O'��t];�SF��L�h���r<���u��|f��wE>���M����
)�3�j�"��,$�g1v��#I���m���"��`6�1g7nh�
7���P*�ag�j:G���}(����c�Y�'1�c)m�yӻ?搿ݓ���|��Ui���C��Y�k��K唢�5sl]m{_���*6��8����m�e�ar�Ѱ�߇��)?,��䛤�a^nI�1G�}+��U�~�+����^���sy��y�{�g��c��d?d�w��y^���6W��h,봔�[��#��>���s������G�t��<��̿,O�t����x���YF�D�����F���vc-���Q����~�����u���������?5sO���3��CJf���]F{�N��]�8���q����O~4X�#s|��|����.�������I���O-�i����Cfz���vciF����]a?e�����t�����Oɭ���=�I��w����@gEiT�����Jͪ�(�Z�9+O�˱��J�R�:iv�M?�Ȱ��2)�_ȣ��,������T��Y��B��H:����g{�H���=�y���"KL9�z�\Ÿ�Ĝ�b|�y�S<��"|ȯ�LR�����/�u��i�ʭ*㷉SX�D�\�H&����"H���|����!-���^z&~����ζ�%��P>�*���U��uP��9mb�O:���
}�T��"&�c�X��� o��T�𪼴%�xu���_��:|.UMn��P�;m��CL�'�t*_}���h�Wՙ!j0��ў��a!��]9Y���k�0���hC�勨��o4<�K
������9�]ȣ��w3��Ì$�����N�Azx�6�	c6���ۀw�P��0�\��X�`�9$�E��
'a��MsX謋bj3�( �[�4m	����5V�Ԑ��Vd;��\(��3$q���O#��a6 ��rQ�A��tw5��d��g�sĹ�������l�|7�=?���&t����l����z�ꍮ�7,�c� [�����$dɎ<�&��6,������<���O�+}BUh�����Xk�"��t_J�~cӁ���9�&岟��FԵ��US?�������G�V�? a�:
����r|�K�Q�s�ہQ�dԵ��A��v�_m���hX/uf���7����F�U�}��9����x�.3�9���3/�
H�#��a�.f1l�f\���M�"�d�xd㐫9���g��<��އ����Μ�k�!F��!G2Mg!'r�V�#0S��x�R*7�8"fC�2uǙMna#5d����o�/��+1��cm��fÜ���Ǥ���wN����k�xi�c��X>\>`~8}��;����A��&)�� �!#�ܨ��Ǎ�a�5��������8�6�A�<"a�Ou�>X���B�s��3i��<Y����h�We��~u���pS�9j��d����u������^"!|�Nm;�hjC�� ���X��O��"z�p�
�!&L?(�����.YK҅u�2�hm_�6�|���k���l�����]@zw��1�bI@�'�.<c���!�= |-����s��;��I��Y�Na��2Yq6�,�:W3[iR��x�*o�v����bg�ܝRC@4 ��v_@��~�t3�̕�(�&uQ�M����% h}b�։�(A7<��M��(�6o�u>J]`�P��p�a0<��ō��R��Gf�T�鰐^sr�+����?�d���gm,��}b+4G���;�k݉�"��������l�\�E $�G�������R�tM̃�,�+G�yl��&��m�}o�1��ƽ7 �x��9]�����CV��&1���u��`2���bC]}�?f�������`�ok�������/}c����jj/V��+9�F��R�M^Uۿ���z��j鶟���j�f��V�!���o�������쫷������A�FF&6��&�g������Ll��RK�����nvcBށ�G���~H&�T	R6h1m`��|E�?�U6��P�:w�_�h����<�WC��9:F���'��	Ei���[BL�WF2ii�L�[��"fxe:ݮ��O��?�`��5Ǥ+���s>��!���1W?$_��9���L.<��D�m�x����X�Y��&aWq�*���R�g�,�J��xc���Ch��Z"�AT�0_oR��KĴ��w˽��j�.��O���A(Z�Ľ9F>3�;�kjA9Y��ɼ��]2���-�ɛ�e��r���J�Ls^X�e�uls���npS �>���O�"����{؄��)���*��Ws(kYx���k9XV��*]G��c�m���Yu���m�[�wQ�ի�ܻ�4%<DJw�[�/�EC�ơ��h��&�S����MU<X���+���Ƌ������}���hʺ�1�&ة��s�Y�d�
e7�8SD��/?+�T
K���
?w�낇11���a���U���¯��A�l�\{;ε!cUx­a�c;<�NO�:	��3�^A��M�T���<d�H΃У�D#�t�h��5J:�j<�5s�u�4���;4+��b����^���ө�ǀt��`: ��A�|Ӝ��9�_\�� �A<�ڛz��B,tqb{L�.f���M�W	g����إ��&l��N���b�S�|��H�k����h����G�KƂy��zu�;\��Gu�Z��{�,�Ag�c��q��G�Β����3Mj���O?�d�������7,��}a��}��U�߈S"�ywΆM/��q{�e�\ǯ֬�ȑ)5O��x��D[�,S
��R��+Dp�B.٨p�F{ �5<��_L��HJ��x��I����}�a-{��]�($V\EƠ���1P�܍�|�
$�����2�ul4�q�{��L�S)0��(����&8�l�����23���f�Ƭ��N׀����{������дF5��X��K���vz�x�d�oq�q8jk�X�ތ�����O�X��k&-L���f�J@�S�.�n|p��.� W�^[3��847����<0v��!և��yXσ��MnƉ�=����z�z�U
ƅ�I4	"YK��T��XU3�
}�a��d��u�M��r�~�˸��Pҭ��L�����|�+�r�R�M�(������61d�T�'�N�s,9j�
��A�ҝoa\���/.� w�d��9r�W��6qP�����Ɠ���T����~�V�������Y,�]��-�؂�oV'�b칵qH��d�'���8ۍr��c���+ �^�����p"�=�<�\�?du���=vf���-?u�{�	���͹�Pm�<�\T�����&�{aA̫�f/$[�O,��nT@|�ǐ��ɗz��2�F�4!�"qTanr��pO;yZp*��SY���鱮p5�Rҭc��igO��1�̫>�D��{3C`��N�<:#^{3�X�c�a��8x���m24�8���bfu�����&�6�m�R$TE��j�Ql��X���"�:��F;ɗ�|��L�t�5��F���j�~��'��7�~�iK��ט�,YM��?l/�X�5�����W_��+L���f��]�k��hZe��(k�fԇVxV�x���}0c�{�}�w<���z-�]x����×k�ސ/�k>0��k�����+��2�O�Y����+|,�ޏ�_$�o�����$������t:��3��N������Z�e�S�举��HɞS���b�ʴ����j���ȏ>�������4�~r��x��K�������_�Y3g�9͚]�f�d�92,z�|��k��������L][U�Y~�1��t����y�3<x՝����7���vɰ�d=��Ky�=���.��ʩ��JE\X**�R�3���n��'B���)Χ�$�8��\Y�e�<,���$[$��F���P6��r�Q=�L� ����@�)nL_Z�Sx[_r̣�����5�]{�B�b4��X��U�X)p�b|�+�����j�l$)��s�}]��D"P���X�����IV�pQ�G,�B�v��0xjyw�.�oW��������n�u7]G=X��Sy8G�ƃ�:>*,T�M_��0�X�H��Pl�
S+�f/�֘|c�S`�*��������z�	Ќ�?�������[n��ݦ?F�y;�ŗ�� ����`{�Z7��kɚ�-�빞�~2�	}3F4(8F����{�0�n\���K ��c&�aO��j���K�L2�����������Q�9��~�#�ZS�F�- �nK�Z�<�hҒ~��46=b9�?���Mz�I���>sg�;��.�6�.�&X@���^uL����%�@��\��`C-
�I�j���(�� �$-�N�9�z�#S�6���hJ�(��A�k����+�*�B�!;aT,��[Iߡ�%�Uc�ӷCdbgrt\G�vs.�Q����0���V�Cc>��S�	// bG'�c!���t�4�c�DL�n�{N�F�]�����3�i:̣�Y+~HX8χ@���ɴ�G3�BU��x��; <f
L@\���Y��J<K,aau�B����f#�d^vs�:�JSv��9c ��Cg5�{S��9��+�S_�kky@��ȧ�F/͍�kn�����L=~t{Ľ=�|�Y�C���!�?��|T���(D.��/����ǗN/wc�`��a4�u��'��)����P~C�?�����,]��ف������O���q\�׮�� �R�.5w�[��]����St��&�ڝ�ݩs�a���+��r����!�ϴ��ϧ��݀9~X�"vO��q]�L�d 6 ��p��Y�*�E��M�y�ǌ�1 ���l;���U�FD��3i�<�0^��E�qr�Kɝ�5��v��H�V�-����0�5F��iG��i�먜!H�=���Ѱ;΄�˘\�dfO����Q�d�x|)����ggA�;�!�o��M)V�H�������i]�yG�O��o������S�F�|1�/1�ņyfe�{��Wzy�|�wp�`��?���o�r�Ǎ��?��_.Ϲ��O�Z��ł�~�<�޼��t��(䓅ֹ��Gl�s�?���l��Gl�|;����k��v��:�	F�_�?���?�+��
6�T���;�� P�=�C՞s�Zͦ���(W�_�_]>_��%�5�|Lφ$���?d缨I�ؤ~�����G�V�CՓMK�;ؽ�*�z>2�b�؋$�7b�E�1��?��̈�D��Cf�ǰ�Rn_��-VWo�B��q�����*	�-蓼��T�ߕѿT��׍%���6.׀sjJ����?Gg3�]���	@��07l0Xia`�W������ę? )>{7+n�#*fj-��EM���S]��Q<��ȫ8����/ޅI���h�g�"C9�/��A�Q��ˉ�E��&Wg��^�1[����zc:t�2D��֝���ݗZu=���ᠢSI��ZU�FY�6�2�3��A�ب>���T/#?	��1-ɛt��g|!똰i9�� 寶�QP�M�\��Lv���>$�ʅABW��~a�_u}�y�z���L!�q�PA�Mn"X~�7P���i�M��^��VJ�2	��PzZ%��r"�WLh%�} �=���Ҡ��K� �U��>�E�Y_$\|ib�6�Dc���rOf��j��DS���b�g?�6���B��T_�$Wm-����^��K���e�sH2�U����T��Q�چ�� k��c/�{9�R�ķoh�����̈j�){�'�;��w�+�`��V"�����w��7��A���N�2}b~�d�D�9��ߋ��{\�cA�#�z�lƴ�;���[�9An��a]g�� ���b�@y��f�*39L/l����G1/�Q`]w�U*ۣb�=���X���0���+$�"�<�n�RG�9:��Ԇ>�Y�T�M�f΍��Jī�����&c$4n�F����ro�T~i���˜�r���7tX���e�ϧ�Is@T��?��d����S��RD\D.�7�:��`��QZ���>��{�j)�w������_�*7G�����ǜF���k�֚2��L�&��	q]sC�PP���E]>���X6�5�\���ॸR�j6��s�[07��$W��uZ�Bx�����K;#�D�#�z�� p]�:F(�,V�J��ײL̛��Q���hu�Šo09]F��A���On�&��e�ʚ���p˘�����	\��j̵��Z�M�������.e��Z���'-��:E�2C���p�r������!+�@g���ò�g(��ib@0`*o{W���(7�]�f���pc��T���B�	�o���؟���n�o���!�MTE����J$����!�����8Y�]w�D0��0��
���<��h�*H�r\��ul[���j���7���R�s��!�C�>��N��P�G�G���ێ�h�c)�o�.E��h8R g���j4^�,*1�1��A�N��R��\ �?�35�>��Ԑ�D�Vâ�t6�O�{:]�e�7�ySP���`Gk�#��L����3�?��L̏Ѝ��t8 �E4�_*�W^��$f|g�R�W{0N�v)z��z̗UT������	��?�%]EJ�����:���i�qB)���~�0��r����b�f���~?�vz�|���Q���w�����?Ot�҅������?LN���Y^�Opֻ���4�P�|���7����7���u��#�%����}	�ҳC�'r��K�!Q�l�n��CvvѨ���&���aSO:O/�O����|��=E�aB�L�>f���ø�Ɍ��2Oj���������r��z������J�d�OL�3�O�|��wz��ǜ���3f��!tTQ���	��J��Pb:�)�a4:L�l��!_�� 3%c1h]&
���6ޯeS�(q`1��lJ�����"3'敹��<E	(���C
T@�GJޖ�V�73jA��^��kŗ>x^�G�4�@�F#�!ŵ�����	\����ن�n�H������l�A��[�C��f��d�g^��ŵ�����W�ju���|��}� ����]/�=C�U�ط�����c�M�s�n\d>AA��dM�b���X�6��Mk���Hz!�:d��pO����ӂ<Х�m�=(�e۠�$�]4 �Q&���$\0(b�ʓX��bF�ElSg�����ڸD��*���]B�9���'|��G��>�MV����k΋F�B�}�l�=GM�;W{�}F.�Wz�^�y�j*Hew�f�r������;`1�!�d���K���4�|���ΐqRL�L_d���=KL���T���r|4���S�?v�+�HO�7�;CX��������<#@,���p.�"�cI��}m��
e���H��-	D�L�<��z� p*\�|�l���5l�3afΠs����ē�I����dc��燳�����B�ze�C��ן�;cü���&����u��I%���|�N�c�0���t�`�sVM�@��YA�:�D!�Ǜ����� VVX%tP��W�X��+c<zRtRT�t_6tZ�\�%M�l�Y[c�}�9��+���F��J���P�Y�c9���{�g�G�ui3�C�j�ׯ�n闵�^a�j��F/�:F57(_j��w�m��D�R�0<Fg�50���xR�:`B�48	�s-�W� ���V�O��}��G����r0'(C����}5�b ���\����c@1`Lۅ��]�V�sE��]{V��
1( �>f+�����z��!�օ< �� 5x��� �-�c���+��PX��AH�]db����3ۗ��`�W|7� �.+����Ħ�M���Ȗ����2ke������<h1���0g::�����I��wj���B����׊�#:�U�!X���vړ�#�͠�- �����Xr�˱[���?V���$3�d�L򁯟(�q�Ď�|Gi�YƯ,�aǼȳ��Kc/.�h$�J:��T��G������!T�?����U�a��ٿ����Ì��X�/��Z������k���=Fj��������ď_�oC�m��X:|0�Iz���Yf�ؐIЇ��_��7;Ī�#�aY��Q��ؑҊ��� ���0oI}���Ojɛb�~/������n���Q2p�x��?ː�O^ːl"Rs4Di��[f.X����l�Z����+d���� �o�����!�dd{���R���K�w�3#3�g��G2��!$����#��E�dc��2�a��j���	y~4���^�!9�e7,LH��r��*u�H�l4�4��<,��oo��܏��})���=�ĉJ����+l�R��$�Jvxi�,��KG~���0g.e�5W�Լ��)Nw��e�2Y�_f�첕h���Mc(S�˙�Gm��E�`�&��t�k4��<�(Ϧbp�[ũS9H�/�C�����Q�w
����K-�:k��Ĺ*�r� ���ddHK��G��Р>�?�||1�k�A%��D��:ؼ��ӛ{�y���å.3AɈu#)�I#"��X��s�>^fE�0?0�ۃmQ{XŴ�:tAhq	��_о���S��+����.0�`C�i})����L@��|���O�.�xM+��%&Yy	��¾\J��Y�!-7����:U�ַq�.- �	*�ژĄ��&�3��Pn��������t_P~�ZY�M'��W�>��D�( �~O�.�M������B@T�T����ҭn����?�E{1��`���{/d-]�HfC�I׫Y%��'�x�E�������X����5 H ��>`]��;f�f�і�� b��&�-���^���}΅��X����\k���v��n����i�7���R(��2ź�u�a��u��_�Hu'CP2X�\�O�4�x�f�K'
�f�c�����gf�y�ڛݬ�8x�g�z�n�_�'��k�`�MHS@��764���@�[S
�,4�kx�o{֖���bPԇ
-3F_���i>���:.?�8p5��ѩ_�N
��۳ù���A�(����� S�Zb`c���d=1!���9q���/-3ܗ� vsI�xru�A0>*�z�D�>��Y�z ���_����Q��	rf
�*
��˯�$�_]Lh������}��
}�S?B�r2Ԛ�w]��a���~j��[��ZԴ�5���9��čbW�:6�xy����A�@�|wm�0�({��}�kq��U,��h�>�+�� ��N@���J�~�"s-d�EʶE�u> �n4
2]���Vp�h\�F<�7��{��\��|�	e��r��!q�������Bq�9H�Q����9���&�BW�s��W�� Y�U��' �(R	�"}�1s}�jڃTƻU��5���E�Y�O�.�I��l� ���9#��H�o�L���;Cz�iƧ�J���_�O\���~���]��ڗo���kS�@{��>!��A%�b~�ct�}x��}.	��G��u�Ѻ�?���G~�7u�S/�Y�Z�m�{�y���t�ع�[z.�4���2�!�xZ_o���<gh�7�族�ү��r�m��o��U�%�^-[g�y_�-�_IZ�{���U��
�\�Y����)�O:�,���ɚ����r�}?�]�'�K�ȿ:��k+���%�PX?X���,���K�n�g9E��x�TX5�	�h�P���_�_n�9�N��Ŕ�؍����+-LPg�tV0񴨁ߨ����J� ��E�v"�*��!��E�v��	:Q{P������=�+�Gf�K��O��bZA�eZ��C�Եq��b��j�{!t�(s��[aU�N	�}��1	��t���]g�z��*��Hn�	 Gm��.~7���Fyo�P�� ����B��<�& u�\v��
+���P+8�����E�J�o���V�Z%���j8��P��o@��mi魰*g��c�عV�M�Lm�\��)�S߀�gs�h�څ�J��hK��b;���X�L�����+������������������Ͼ���˓{���Z�^��V��{�X�W8uw��P�-��r[�yeK�&}<�Z҇�
��NY�İ3f��@�IPS���{,��(���U~7D��o���Փ*��u��E�GS����0^m|"(�!�����nʳ)�U"&�G�Ou4�_B[�(��~3��x6��0O�kG�?�&pB9&�F#�G *�#8��#�f�d��t!ʃx�$F,t�^�Q_y��χi����#�� �Bh����o
�LW�쯀��7{(�~]]7�J7�.�vg�v�5��`��˘�	�� ��w��=��y5�	Z��#�k�{�ŜW"�!��[�Q6~`�.W�W�n�O���j���^��Z��n Z����4_o�d��G��l���uu��b	C���p���y��{Qt���ck��}�ީߩ�_,��R��U�E�\@�ٵ�X�p���pm�3KS�eb�:ڽ?���C������
[�gR�z��Ʋ�
X�
}?md��������F�^n��+[��e��Ā�B�T~c*Ϲ��""S���Q�|��=�gڃAgK�ۃh�=���),���#B-?�ˎf�;���lޫq��1I@�D��`�羷�o�����&Է^��|���s��0��G�����D��S�*/$�]�9?��┡�0Ѐ��S(����Ř�*ҍ��և-S;u�p�\훇�h*�$睡Y���qbP@#�s[����t�P����!V0��ɓ8���X��v6s̳I+8��݉?���۪�S��?��w���[A-�������H��4�b���?*����o��T����J�S�ָ�5�b]Y|{�mY��ߍo�j����Z�}$����e�����,�OU�ݖ����_����������`�Ơ��^������]������_�O��[���E�5ڟ�z�k�:�����;�ݿ)�O��������� �~��6�����j�Y��_v��\�1����y��J�ع�>������ם��ř��s�I��\z�,��=םw����d��3qDǻ��|�#(ߪ.�ga �)Ȏ�b5��R7��=O �1G��3|W��������j��P�ū,�?��ȡ'��e��+�mY�ʗa����J�������,,Mk�X,�Wb���Uz����7R�o��"/\��h��̓�|^C԰VNc!��)g�q����j=qx�wǪ��:��g����ź�n�!(�݀�?j�x_(���2�Z�S����(Ҕ�Nݏ��ĒVؕo�e�U�b�N�;��Ju�]��8u�@X
��/�z܊.R���24ٱns�p9j�:�mBb,��#Z��	M;���h�YE�s�
V�1a�����}B��3��d��1�+���o�(q��R{�(�&�S9�}p�V)�Z
6�6~��t>yT�`����m��~�03dsc�����I�������Ds�#>��G�w�����0����8���*ڈ�p�����F�_	~�tR6Uv4lm2���-�b���9��9�D�Z_ճ|���b
���&�$(�p[r�&�G#ĲϰK��a�|>l���N�Y�`.0�����U fԘ�L]�"� �+�D2�:j�8;t֘2���q��ڎ�h:T(q\���2E|+D5xn3�7�:󠗙�S=s�������Pw��_���q�N�OX�̵�U�>_;�|��U�lU�f�����I�]1��U� �=�׺�Д#��
��b�5qZ��õ_��k�mS������,2���uktP�D)��}#��PVd��i�~��l��]���J�!K1!
���[�s���(�tx�/�D;b��ѝo��kb,�3Z	Q����LDT@\��xZ�[�����fo�&	�:�B��(PŪ�"�����!��SX#Ǭ�ܢ=qQa(��T�t+k���92�?���f^�]�"$��T>��xT��IÓ��x��	�)�,W�*E˅b����/Ç�~�P�^#��c���v��U��F�|*E���+����w{�%�|1�=gX�ym��ƾ`���y�+��&۞�%�=��W9��~η)a��m�����R��'^���l��QfM�TF*V�ugE^���3�_�e�cv����5���ڎ��G���P�i�����8Y�8���^c���g_ȟim��,*Y��_m���D�������/g+.&� �R�ԓ�u[y�]@������Q���Tv�J8���_t^]�����A�O��E��Z�%�?�c��r�s%��7�f�����%-�a�j��.�8�w��p�= �k�T榴��K,���/��e�p6�+ד6��}��}0y�U%`��z+s	��oPV��J:_�
�*�S��!Vķ2�	x�6MPմ�:Y]g�����e!Z?N�/��fm� �i,��I*卛D�D���Q�7�7����̣�o�0󃾡�n�_��:ãҮ@@����؝
��J�U@��*�X��ݼ�!a�*�r/�Ǣ�m��ΆB����R`X�Hե�3U�Mr�ۄZ|�g��i����Ѷi_m[C�V�߶B����~�}Ա�*X�U!��e�J���SU*a*�Rw��P|1�\yd7����Rڪ�b*�N�G�5g��I�Q^���>�ܣ�c�9}iS#��j�/q�4v-$�1?B'����h��ڔӣ�9�񸿑�Ә��E=i��~�	�Ye"%���h�*.f|,(4��F�g�qZv���hpF�Z��Lat5�׋7C'��E���0A�n<JnjGo{\"P�����b�c���Sҍ�v��$�oL�}t��a�kcщ^��|]��h�&��=q�����A�|=�0Cǭ,�|"&d^>P"{���T)��Z��)�	��_�( Ċ�}�Z)>2C��خ�������ڈv�]sP�����:��	�> T��벭ު%"Jr���v	�'q��σ|�B����[R,��X&��/�F�0�u�IP��V�7K�[�����c5"SVc�zSu�����JՒ���ր��Gh��$-/�AB:8qP_Ӻ�T�N�&ސjc��S�u�_�	�:t�=��y|ڒȾ��{���tW��v����?9j�v���3��a�FV�vc���"���%�I���s��Y�[D�D�A���9�Cl�?|QY��������J��$�)MT�b](��/>�O�s����6����:�`#:�������rQ�X����	���\����%Z8�@�;qah��7�%ӡ�ij��Q�my��,�*�������H�.�����QuY�,����FuVm�gSt�_��1��<��(�J����aɱ�w���)}�O��]J~b=��"�_q����K�d_���?�W�l��T�d�75��!q���XV�Z��K���_}����\0k��gT��0[��t�"hr�������\�=�N����(����s(G�Oc��:����T�O.�Β3Jדmd�������t3�]s�4f�<���=sq���3*%_B�% ��ټ�Wug cz����&�R4,YN\I��1p��M|����(-b*r�W���puٸո��꺘1s6�Q�2���A/4�ѥ�yT@��cB��F�U$q�?�q�N�
ՃZ�>� �X�
�XZ���搵�.��-�J�HD��.O�ͻ��<���*�u(�h�~w,E�\N�nBH��]]O�v�����.����+i�yx�G׃mU�D���#<,�o��:"B��>e�Q�{6ճa�:�|���@L(f��~+���*���~��^�%%�~�h1�hX�5 �u�d����lg�vk�37uW?�6�|wS?C^�`��{u����@�	z�3s*�ԛ1�j�]��J���a���%�:79��d�h�F����y��[��u����[��o b�:�ӛ�@}s���(@vr��&	k�OZt�x믣��.|ޮ�>?h��q���r��W�(�!���t��o	������h����q�#����;���`�rW{�ȹ��a㌎�����W��/b��4d���=.6a�ƚ~�S>6��Q̔@q����=�d�{��0����WWH��|"f��otA��*UE�W��Ϧ-�
���e)k$:Ύu����i+��p��K̾�眸���#��+��(ᭂ��b�3�F�d�ˍ�%�&���-uz��
�q�V�Jޚ���G�y����RFcmuy��R��:Pvf�wz�D�FC�	�Ś�7KM���FGc!q[v;[�;'GQX�5#�A�9�����XQ��S݅��m0�Mx�ñ�&��%S��+B�Q����s�¹�𷲔/����ǎV�W�؜�P3 ��$gn�ƫ�h�c�����}�b"�d_���B�.��h�ҪGs�gQz0k��C8�P*��:�b=�ix�δ�tB�Og�}:��a�\8���wQJ�Yp!o$��m�F=G�����糿�BT7k��l#)�z��w*����1��	;��9/K�c���`y�R_�iuX������?����V�>�o��`���y>%5�lwlX�k~V��_�;K`�x}�`������k��ĳ�V�$��r}D|�q~�5\��
?��9�O���~����G�������fY�Uޚ���Ux5���z+��^�Я��,���_I*_��8�q2�Tv,�uO�U�%�}EOv2�}g�E��Z��+[����ڹ`��k�i����%�䧱��_�H�,��
���z��a)�{��Q�u�j�[eU����rL��w�7"�j�4���-Rhq���AD15>&�y)z!�u���_S@�+'�L���ug��t�,vI�A�e�7X��k���"2����g��x3�:fX��1��Tر��&WS������6�? �J5��T�7YGթqjU��u��������V|�F�{)"!�
����z����V���r.xi��8�Ő�M�[�̼�h�����*L���T���I�*���长������tv�+��Be憖ehp�}X�ZdvC��f��_\3:������@�PC�1Ul����\��X(���A�����``|'rY�Y��"�z���it-��g��Վ-a�C���uxW�R�}�nu�wԮ�q�ч�i�ߴ�+w!�V+��:�Z���}S����ĭ�qjzn��6�`t!�]��K��厇 �xA��F�\YJ�0C��$��W���0�^nԆ��R%3��5D�Cc�a��
�f͟��&��q�;��p��;"��<_F07jF49�[C�Hv�F��"Φ��Pb���͂��,�Ta�7?��P��&��=޵&u���ʲU�|�?�6<N��)��y��Ԝ��e1P��E�Zʖŭ��۵���!7~��Y��]�PC\5�s]/sQ�bzw!Q�KVD&����
q荻����L�Wt��qa��<*��uu�7��H��0�nZ��t�Q��ky-_ǂ�v͕���%~G�_L�&&����`�r��r��D�6�Jw
�бL��0���8��b�����ȋk���%dgfU��m�{�����5�.m��*6����D�M��B�Ř�u�������ApU�b�#4�o�сA��u:~���QNc������������O��s#���"������4/�ŭ��d��ȹЋ�a�s����� �(�7�<�����[�1#��n�en9-?Ս��9�P����YF��cM�b賞��ci�>��O���~�>�.���+�{��ά/]"��(6���8��C�5�o���{L�z���ޢS-_������K�zYK�O��U���9
��'��
W�N�����ժ~���;�+��^�Ov������2K�>*�_�+��6��j+�d��� {������s%h�����������9H���x�'�B�U��mN\.g�Ι+w1�L}͜��X�[���~#c�U��|̙YxV�=D���Ƶ�D̵����X*]ai��c�S���Ɓ���֑�s-�"i�t��1��it��$�Mk����[1�?\p��&R"�]o�{�����Pz�n���.��� �"A�fd1� ��1����J�t����bŎ�H�XSǻΫ����DbF���p�̯�虺�ϩ���(�>���<��z����z�=b�N3�(���.J:Oۇ���ʝa���D3��C��&-^l~^m�̽m�P܊E���	�G-�o��Zz(.��c��Rw�R7T¶���m*�y�<,�c�@�%VH���߬t�
��ṇpG�F5�1��=S��Q�iy��*֩�Х�Φb@��P,v�-��o�j�{���d���>�^�-�l���Y$ �J�'��5�Z��i��'yq<���O<�2�*�o�aa�/ j��d��
A�6c�K�V�7�N(O�F���HD������CR:���>:쟀����h��	�`E�5��OU&јXE�h���srQ`��/�ݸ�Mh����p�8��p�����îL@�[�[j��D��Oa����4�߭d�K�����֖;���#�?\���T+5�u�C��\� ��&��9Y�\9T>��l��������`�&�2^?�����?�,���iyo0>��uLm��S�f��!�I���&��B�9�p�k-7��0�k����y@Tf:���U��Thu��h�Ԃ:Ś�}�^'��-Y�y�Y�!e4k�!G��ږ�6�ε���E1� �����l9�#
F�1uȃ�.'dqk�>gz5YT�X���'s���&�јv�.mw��be���6�{����"��4�=���93�$�+ȴ�e�_� ��|�����p��~:Քb�W!v�F��E%|��E���Ly�R���a_�k�G��A���g��T�f>~�~\�~]�Y�a�n�M��-預9n ��e�zס�~�<�p��bt~��S
�}�+�m)h�{���}��*�qj����<dPYܿ�=��>҅O�H�žR������Str��4,����������\�n��~s���6r�� G*YSZ.F��=�j�e�6�'\���)s\�hBFv��Q���W��忾�	�O�%K��l7�۹o��F����fA��wH���(�M����j!^l����{it"��5�����X�5�|�_�~�!�l&A���Y���&��4$	�8y�8��Mn���.w�;��@��6����^�&sՋ*&�8�urBB�3*�7�Ζg�і�΍��"C�.�s�;%��6�kw��e#%�<�NY��g��l��N�ga���X?�pͯ&���tǄ#��V�5�{�=������~��ء�H�3Ϸ-vZc�y�b5#>bSn� O1�F����4��Z�J�)PӸ�7��b{��S!@��kR�Щ{c۫7��C�r*�0]g@�ۄ1�¨�$�;d0T�����W�i��Z�do���,;����X����N5�/#}�:.h�.���Z�mQ7*l��0w�-��#.�+��-���~?̀��'�x��2�H+�h�d U*ҩǘ��z�8JEͤ��ѐ�1)�D�b�03�Ԗ�an,��j�(��l"J���e�Ӧ���+� ����^c�q�����.f���'
��W�j��Z���:�V¹X���,�hP�g|������2�f'�!:4n{RÞ���b�qn���ѹ�'���F�w��Y��^(�9k�f�롏^��@�L�|�����ֽe���J�����d�;V��,'�?7���lK$���Vë�]1*�������8��?��N~���?���Z�W/F��b�o:/Q��!P��:t��_���XBv���C��㾫po#���� �3�������N���{P���a�~��]�N�Ƚ�f���d�d�͚�z���A[���-�j߭�U�w�!���Q=�Gbċ��3�9��C�#��z��H�As�+yZ���YƉ�`�'��
N�,Cxu5�����fd��,-=��G���)�ڹ������}��}�������7���/�ו�Y�%�X`�u�S�o���yך8|�b�����/��/���/�xI�_b�ש�],�d�K+���doXڗR�%+��9��]�Xu��W>7�����Ƒ6�l�UGF�������T#���L���;|�=�,�o!�1��b���׬7�#ȟ����?����FP�q���Z��>�׃�%�bI���7(�$�X+�Y4y	h)+K�E�(��L��I���⾺d���c�Y:V�ePA��:�>t�0��G
i�B�^l>�ɢe-����'��8dS���f��J0��쿄JD���WC� ��2��j�q*�F�uo/	�ܙ~�WX�Fut�������8޸zC=�\|�j-�[d�l�F�O���z������azq�*Xkt�qV竿\Y�~�q�箢��nvb3;�b}�DCK�JW�Imش�%T���=K�Ư.�A������Ʒ3�-,�o�F	q6q;G#�8sp������%@�3�(�ryݟ�,�"io�����ޙ�]wݧ��R�n�?���J�&;S��\�r����莳Wa�t�(Ȟ������̅��ɸU?p%��&�?DA�d�
�_,��>x���Ё�*���*L3֍���hD��?���Fv�]b(��1�r�����o�a���p�vS�Q�}��������@v<U�fz=6��z��%�c�c��7�%gW�dƫ��(��vԐ�	�����* f�`r�3L�j��]t^s�x�^I�鐎��>q��W��mUކf�ߦ��jB+2��R^�ym��6���K����i{�/����A��ߥ� �]J� 2cIW,�!��AQ���U1��Gf�J[��(�Wc�K��4��j�v�v�B�h܀�cu�.�Ȅ����B Ms��@����-���]�j(������x/:�[�<j<q�~j� ��Z�G���"h����Ge���ݸ��}&�-�������
'+������=��Y�Q2�sl���&�~Gҏ�>����]�ʡy�{��5��g����a.�f�Rb[�o��&�1�?��t���\£j0��U�K5?�wh�$ ��Y�8<�ck�co4�g3f��}� 셱M� ���"�W� �I�̿��[_��+����$D�2j�"����%]|���������5�������$^��w���g�/z�b����1"/w�o�SM����Rs�|�9ž�̉�+���(?fIY-If��W��-�_��k�̝�JK�Y��ke�����g��!ߩC�\_��kN�_�� �h�}-��C�;�Xt�)z��L�E[�
�6�%������5b���M,�S).�W��.�����1H�*�6���H��؈%D_1K��S�lҪn�X����!]�����Xq}���C�X��wA�X���K������!�T��ꥶ'�T��l����j�QVP�V)�U+����	}Tb	�'Myb��?�k���o�4&Y���ݱ�y�Ѹ���怶���>�i�"�h�@�
,���F�� ䷷��JQ��h/��;έ��Q�2G���dM��15��~�:)!;Y�gښyx-:J��/B���1�(WD˫��1#�ץUHS���	�\KdI<|9]��^�hwA�^�V]#y�NR��@zÉ�73.��1iE�}G��� 8�ӏEw���� s0�		�&��ݛ�pB�%駿��c$~~��&!`wv�Rc���
W�.�
��ʏ0����3ǃ����u�o����8�T�L��G��Piܜ���t~�Q3�m��C�A��Lc������.�y��cO�ױQa7 �q�fm�������=�a�g�^� ��F,A�K
ȸ����GQ� u�P0�p6G
q�2���~~)���F��~���:���?o�t^B�z��5�*�7�i��t._,�Pk��]��\�_hUL����(jA��HK������XV�nE�i����K���r�{�R^���_�_K�)�NVV,���R���W��|���ˣs�2��qp|���7�]�v��lW�FQ`��n�D��}��?�����/�ϒIM�4e{Lf7r�n�c��˗��@GZ��N[��3Ѕ��O�}6ڗ/���@G���c�H/�����MA��=�/����&��I�E��!�谈b	K�h<�:���@�*��Jcm�~����=�M��L��=t�ϻ{|i&��w�����?�L5��Η��w������o�~F_��wT0z��mɿ��_�ȗ���/��w���p>���+��e������c|Q^r���~���7q�	���1{ �P��zS	;�&!�Q!�I�kh�F&d�g"�g7�/kӏ!O%��i�7@��g ?=Ǎ��ِ>+������.�^m@��+R�)��������|y/�ڸ�F�S:nQE"v�ƭ
�2'�	�[&=IY����p�����G{��p'6J܉�R�g�Q���Y'썷������{�v��B�֑4E���q&�%4�����p'��W��`_�q7�;���T��;�<�ؘ�!_T�w	���纟�G�$o�����!Bb+�8�бĨ�lP٨78!ñ������(6۳�O{���[!���h�԰�2:s�v�D�r��:�YM�k���4�뇔�p��m���q��Tռ�)�"ȹ-2"��M����[icݴ��:<���kR�7f/p�zť���6/iX� ��Ƒy��|]����C|_&.p���=B�Ұ�	�O���W_`D��M��!=�HIm�.��]�[D;�����M^A��7���C����ȼD��(�Tӑ�į�K\�.i5�&�R>(�σ�o0��0��0�{ d�%& ��1������, ����ildk��x�D�鐾��o�@�q��S	�,��N�^�	0�L���O75��Ώ{,V]ўܑC~U�B0��g���'���?�����_���$��	f7L��.��%�65�t���L�e�MP�ъ�Լ3�c��a�65���F�K�� ���U��V%&cUL�{�ĉ��(������n$B�1t��������X��F:��
��@�0�X�Qq��;����x��a�9�d�%(^�A�Tq�����U�w�^���@>j�Ny�T�8�I#�o�36=跢���h�F���l� �B�p�V��C��>��΃��Q|t�ι��L.�WZ�S%�7n�Ө:���X�]�Е�l�����u,1M�X7�N*���	X\�Lrb�9�^�g��1�xB�KLLB�ƒ����a�l��ך?�M;�K[~����+��%~���/E�ŸY{e0�k���L��(4���_�^K��?�fR_��_k˵c.v}7�w��T��˾�����{io��@М%�kx���}�X��d_��� �}��-������?�������������l�_^8��?�#.�8�^3[z����^�<����g%�n�V^�㻒�c����>�LY��[��#6�kGĘ�
�Tll��p�Ȟ�y��?������j/�b�L��T���R�}�/����:�����xN�����,��-K-���j*�S���jvS>�
8�a����a�:��b�%` W�&��c�S'�����TY����ϸ�
���t�h��zH|�i���~����GS�G���@Յ�H+x@7�бDp+ߕ�޸���}D���a�h�%�/��]7 ;��W��-kk��/��/����*��\_b	aE���!&�_����R� �~@���
�?br�,�K�-���̗W����������/O����l��`jb����`HK�\�R�[�ț�`Z��f��7-��xΰ�Z�G��J� �;_��u����}������@^=�����u;��8���q?H�ƭ����{T��7�.��-̔:^���Y2e �������r�cN�+�EOz��n�0c8��F
�1���
3o��j69�[4��!��R����d��!�|0��_�	$�	�?'��$���X�`?7fp���)? �u�І�p�t2�Z��Y��q��*���Q�.�܉f_�@T��C8>���Kϒ�f�ڿZ�}צRX�g
��R ��t�"��&�B�p���?�̶�"��v��[�F��n���!Z�M�&�[�����ė
T��}�}w��|a�FJ�I�j�gm����{mԵ�ށE>Ķ(Wq�?(��aļ��0D�5A}P��¡s
҄c����TD�w�k����L��e��*h�� B+��^}rZ�,�ę�L��G���J69���o�z|��������^��}9��d����5 �ZX-��������y}1��a�ly%<_`�ɸ_�_`��G��_~�ZY\K+�����~��_�p~����?�B����]oC>�5&�9�ޮ�]�o|���θ�g���0��+#����N�>Ptv㯯��'�6C����ˏ����!���fN����{��!9��w(�Y��zN�,�h��_u�j���2�?6�������=d������ۘ� ���R6�t��_�꣒73�jd���k��dD�c�R����K_ǆu^,����1/�3��_��:4��s?ñ�A�a�y��Y��^0�:�:��Z�cI7��k}�<�n��P�T��O7r��t���.w��r�)�i��*}�9ؤW�I���>�h L7��֑ٶq!����Ԯ�4���I$I,q��I����߱xѢ�_VpL�=�, =&��+�5�V�7$7�qh����oܘ�q�E�m�l�Ż�± ��o�㜢гc3���T7a�_�Ѵt@n-����h�N��]���7OB�����Q�����S;��+$g���̒ثġ��P�;���$,��|���b4Tw��3�X�7�4_��.�w)ʐ�lO5۳�Y��d�}�Q���ɗ3%hFmk�(���|1Y�dP��y�&
�����g;�v>�����S΃%�=�3��0 �Ɋq|(j�+�bX��u�^:��Wd�c4b�W�\wu#E;f��xϝ��&������&3�?7�<|�ĥ.�����A:^��C��U��Ѡ��҄y`���]*�n�ynW�Xǭ��^;W9�ߨH�𣿆x|���@��l��N��7��X{3O�K�����(2���8E��~1��W� '�T0����S9t�H<��8�����5���Bp��܉�:��/g"�ǅ�N0|����=�L����E���<gO�U)t�-�Z���4���q���LO��C>K��Y��>/(��0�͇���A֭b�m��-1�w�����1އ狘[�?�ˀ���x�|/���u��B}���5������w�M��wagg�R�"��;�C�͈旊��,�����?���ߧ����5��[��;;�����x���/{����]�Wͮ��5Wx3Q�y���=�y|Ph�+��6��:=�:�eT}���Ion����E�K(cI�w1��z��%bOJ�(���|�|��^��O
r.m�pM�:�L��������6��&D��z�y+�5��?��?����(ȷj!ְV<[n�(V"�b)��0K�+�:�^� �Q-�~�.�$���5�ד��t=���s5�
4�V���8v�0/�`f��F5�a��d���l��sZ��^�q�7hM�|�/����A�8(��{u'�U��(�7�x�	I=H�>��y�s��R���	�m�+)Z>�Qz�&�� �Y�ݷ�x�����9�%�b@V�>Q2���b?�Ǯ*�S$��Oc�ǣ��C��u��\����;x]��/��#z�*x�Qi"�Q�#�t�"���-� l�b)﫣�l_�,��K��}t�X@���X��z �(%x(�I,밞�V\)`���q�ŷj�]|Dn�`;����3-4��PYE!���Ӂ�`�� ڸ�s&�,U�5�,�%��
�|~	��:����*�2��6�Q���S�y��M��hh�.�NE��a�jh=%��\�xe�Β�
4��ΫpF���M�Um,�@z���iiP�/]�n�.���յ}�� �Ҏ�`t�+��7�1�}m�S�N��Gge#�:���U�r[��1«�,����u�O����)u�.�7#��βD4{T�|_Duk	s�T8(�BtE��,��$�B|qYX/WBx���i���83�2g;�g"`;n�Y���Yj���و�φ���Eo���o�����m\�����+�����Ï�u}gV)��ݷ�2�V�Cv�3�/�W���|'/�s�~� ���o!s(B�Z��g.f}/�M|���>;���F��̆l3g��U�c&�y��e����<0�7��r�_͚y���H�~�.f�zm��d��{n�JE�u̓3��`��f _�r��eK�s�6ZlW���:��|�\�#K�'��,?�x���#���Kr� ����K�T� w�n���
�?��|_;����n&  D�(gp�����"�;u"�����.��x��w�T=uc�K�n�u��&ᇛ �z*�����q{*ޱ�L˨.X���
��Vԯ�;�J_�[:_j�\}��86�>q[Brl3��`�B�i]�f_|��D�&q���ĭ`6{t;>��ݟ�Ql1��[	1��P4� �lͼ4������T��1��>:}n�e��E��u���(��n�i����5V��1�׺G琿h����׭62x���y5=���W�AoT�2�"�i�3Nn�;� wa���=!�^+"�u��>��ǔ;a�DǷ:�_�Q@1�@�ϔa��V߆[!�G8:6�!�$� ��������ja)o|ӝ���q`P3��!k�l㒻�I�B���1�e�g�P+��JކfC�1�s�6�l��T��9���1�=� ��ly���%>�$�!���{m*/��,��;>GJ��X˪`��>�+O�K ë���4�L����rN3�J~jc��QQ�ZS�#�X�j�7��߆�����*|��w!>�Bl[��\}2G%���*�Y����a�vl!�6��lm� �T�?�i�V�K3���;��j/8=w)_�BH���;?Z��0��A����}$9>*�̟����_Ʌ;��6ï�r:C�(�`��'�rg<�w?�Z�Z��F���qUٟ��Ł��y�Dem�ZxN�W{�����>/��[z�T�����AϬ�����`[���v=k� �/�T�hă�n�w�U=|�Ľ���A�J;~!��N��Ȝ����p�lΓy�Q�d���m�AR�_�N�\�����z|VK�2ajΒ�֢��*5��w3_�z�+#�����!���}͊�Vz6��� �053+Tem�d��h�ԝ?8��Vq�\�Dҏ��n�L`�2������0)Yݘ��[7�%��!����xU#��V[�q/:����W��w�@��w7Ɯ��/Վg^�o8�jW�:����>�	rKrh����K�����7TM-a�PK@yq�d|�n�yi�-�3���
b�
��%��?��W{��j�^�^&^X�D�Xo�}��9j_�;��� ��{�o�����n��+k�IuAm=��7�A�ޤ�t=c)�� ���:;/5\3K˛B<g௭eh=�	KQ�����z�o�5K����^��/gbvK`��歶��﵄Q������%\lc	,����؆ [�� ��p������GEa8*s��){S!=O�53���*���*���}���ؤU�M�F,�6 m������)z
P"O.�CyF���b	��C,ȭv�+;J�
$O����e��gE8[���Pߩ���XE��oۈ/��%<���ϻI�&J��-��t��.���h1�)������x�W�/,A]�g(��|�ǳ��Lˣ|��){���I^ڤ_m-E7e���[JL�bu䋎�n��f�%"ޮ�a��
*�]��uF7�b���(ڕ�=�.�0q�X�l<V���o߱s�G(CS��C[�ҠJ��:��8�K���a�
\��i_ 2��y�T�­)�>h��������<TC7,,kYz�+�D2T�[=�����,�M�K?JK��ʤ�4�FNg"z�T����w�&QX!��Ī����yAG��ZY�2g�VK�ٽ�^W���)h����E*��D_k�ȟ%�����/��S�|M+�W�uշ��"��:���V^�/<�^z�����yA�Y�YO�A6�b<�R������ן������=�������'��|]����I��������>	�3+��k���	��-���7��9͸�h��Jo�[�o{���]�b������W	��ԕò�����Z*����d��n�B� ��(i��� @,6���/��|�R\3�ّ���>�NT.��e��N�M����?���!��C�N��R�f�=�j��r_�L�Ê�k��Ю��X��j���������\$��(0h�k�&�;q窳���8D��v�q�UJ|7��`� �^8�G��������Ky끋W��9Tf�Ek3�� ���χ �V��W<����MP��#�|3��@>�r� ���<�l��B�]�b��{t���{��ʼ{m^�;Q���C���|]���X���~pc�������t��u#(b���:�����8_�Dt�7��~��:�N�ƛ������s!�'�:�Pe�p��q����Yю��~t �Xҫt �v��[da&ʀk\b_^��z��yI<�F����holT��2�/[R�ѸU���\�r��$��y��ҵ�HK���^�P3��U������Í�s���*�;���8rcK�����T����:Om���A�Z�Ҋ�*czbAk��7�a��ȯ����;������NK��t�]���h�HՉ��%�)��f����S#'Bg�f����nP;v�9�x�ݱ�؝��ְ~��.�$J�='��Hߺ�?DE\Y���R/�Ak�z,�m(N9P�Jwr��=���(����x<CǎD��Aq��S���.h5qlgj�Y��\�J�*.u�%���-(6~��,�^�x�J�+��+q�p-��7�b!��^����k��L��#��������|������ZEܭ�/�'����#�Pm�1�l�1~M�VN6Q�]�e��, �#Swˡ4�g��=���,�f�����H�;b��FN�P@��Ƭ�.��M��~O��w)�b'��F܉�ׄYQV�0�6�~��7�X2����i�5PkB�q�-p^d��V�'�G�E�iT�r^:ڊ���D�	�5��\�NDׄ�Ա�tfEN=��\��"�<�+��[<mo���H���.��6_|���m�Z��U��Շ�,�*C�(��yibM{�X���n�"<���6�m��֜ �Tzc^`n�x�����1!m�@l�q�vIy�A��?�?L3�؞%�ݒy��W��g	�k��uŅ���e2�Yڹ6��z7+v!p+����1����䋸�wiIu�e�b�`����6��Rߝ_h�@w����1�����+��18���@�Z$Ȉ�G��F�%ޫ�<[M�vkz=����5�ײiv%�}��I�zU��,�;$��Mh8w�c(��?�1��<cd�"U�ϻRs��X��Jf��du�>4���D��w�%��9 ���V;',�9Ak�)�1/ x��M6��A~�qL���$�gh=[E���SɌ)Ж�ȸx ��Io�n���Qa�w>��ص�&�*��R'��;J���zTE#�Y��5v�X�FK
������q����v�_*:l��ilBP�
�ݵ����z;	���0�5����3p|��ĔقCޤ �9/�N��2�}�\��#$;�j3F����.,�0�ҁ�:s1�5p]=$qwh�˷�?<֪��6fky���1��������W��﷪�B�~ x��2���\�wmK���A1���/���|�/�m�����}���y��T�.|Xc��`r�7U����
��3K���mf�=���k ��r�w��x���3�qoe�HF+�\��ĖfsCR�	&]$���&�R^T��Wf�Mä��"-��Q�8U������-�@.�t�jJy���S�q���W(&o�����L�%D�rh\�=D%�[��@���m^P�=�$k����],������*p�.-I�=��T(�
��U���I�8f�h�� �&�@C�lk^�qt��#/����N��Jمw]��7@���?�/�(������i)���^S7T�.�χ�[�99�V{}��M�����x%��qr��i��$t�O��;����� ���%��L�)J�P�(H�F1���saF<�~��:y�Q2 �b>�O=�9���Zț/JS�(�hl�&����zv�t2g����q(1�a7���YK��YA
�v��a	��4=�rB3$�ٶgGBK�A���wxU�S�{"��M��s��G/o�s�fpi\��_C\Hy�w��l��&� @��7��y�ty��# jq�)�����KB�^�8�� �8�V'}auܹ��yU�i8ܡ�_�!�Z�h\�8�S�����&rd ��\�m���ҹ;W��l,�r��@�:=��� ���=y�-}�6�Il�и��>�o�ӹ��cv���H�}�_>��W1���Z�!��:�(.�A=���L������@�3�y��8:N^�*$�x��͊��g�<� ����v����a����ʱ�~�ε�N�eg�o��}��e��W$��]�����g�w�eb�a@��C�"��f즽F�++�`�����ie�܉8��k��*�2�&qcZ������*l��j�K�_:��u���m�����-z��^{�b�P���#< ����<�Jj�$�7�!/�<뎻qZá-z�\MV�kǼ��J^���%M~�jv�@[���&�^r^bK�B�tt:v{��Z�Ӿ��h7W8-U��frGk\�0��V���5��o�Q���}i���w��0��Q8�_��	UH/����'�:�6Lu�M�,���/܄̾�N�pTڐV:�u}��@���X����%���Ɓ:��0zT��d�9�*$3�9
f`��a�����ܨ�20 �R�ӱ�e mTδ�0������%��o��A��c
'ƨ���U��m���������&WcB2`d.��%�����(Ր�!ʜe��H�o��ԆvdvҺ�ʪi^�:�M&7z6cE��g�OG�'�g�p��q.v��0����C(���^>Hq�B�)d��x]���+�-�Ҋ��%L�*2��PW�HY��/k($���%H��c��&��+��
vlk�4��i��PpI+�X�6[�X>:x���7�� `��%b��2�g�:��MrHl�$l���_�v��N7�7��S��	��2��{m����A�,��j=�r���[�(��Z8��U����:#>;��X�E��3����@�p��d��I^ř*�&l�3�ܯCE���f��C�t<.�w�Kb#Ր�R`(�p�/C�/���u�#Ֆ����G�]�^_k���]O���o���1��S6r�������(�2�Q^7׏M&��4�4����y�F-���έf�Y�3]s�ye���)B����&+|bI�����̴��>��<T�O��B�?+(�*����U�(���U
f:���TpJ��:�H�m;-)ʿT#�wy��1a���2�*���U�瞦,ءQВX��@�K�0���8F��^��2�Z�M���Pnᐱ�zP�5�c	.З#�g�:�N�_�Kޠ�$$��El�yMޏ�5A������̵͡N�n�L�B8x��?4u��I���*���b�����ͦ�B,!����[�
0�	�[@GX�]J7�N������@�2v�����w��W��A=�5W��f�3�~���̉K��!��U$%�@ZE{	�d���t*�kf,��}Qs���{�C]��O���J�%(����d<8E��Ԩ���U��(�D�ȯ'� �5?�}�[rt��a�M:� ���!Of�e}�;�<ac��I�w���=d��)����8�;a�5*�Y����+#�W�&�
��*3����.�&�qjs<Gˏ՜��S]��a��$��)�ƹ �~ ���:g����qt4���f.���C�M�ˈR��n�U�#�Q��r����~�Ð���x�U&S��X��G�o����<��3�C,�{uMĞk2�Z����&[��%��6уk���:�p�����Z�d`���3�֠��k7�;�Do6~e�=��]�o�/K0�&{���M�y Ia�3��~CqV�M�A��C�
��S!uD��zg'�-ր x-�������MK����>ǰ����w��m�.�� �^ �K' W߁��Zu��cu�aY[����W���'��+����J�ب^ߨ�����z�G!��W/��o���-��
���F�Q�f����FB�ź�}g��&ŧ���*��	Eܯ-���*���3}�-��|��:�9Q=����U-z�jJ�	\�})�^IK����fZ:���C�C�\�t^Ң��M�w)��\~]Q4t��V�Z�bԺU�a�y���RמjL,�'��	�u1/����n-ڷ=S_n����L��X<\W��I���hhJ��y����	kS[��H��;�4tSx�f+��d��zSi���A@�W���R�X�T��޸�ް�'�S��D��'��>I)��r�`um���Q(_מƤ���eh�x�2�А���vt��nBHjL�1�b�]�Մ�e�s�����jl�چ����F�!�B �"R�G/�Ĩ0aʔ��W�K�l��t玾��?�#Cy��Мl�3�4TU$��]��dA���K���|�i�Cx�*l���yi�*��4����	u�&��� _�n6_�=�g���M N��������T�u���d�mx[w��g^��ԟ��©�rNw���<����v�K�;��U��Ӕ��H�P{Iػ�y>j�p��K�c�M���(�/z��R���ٔ�m�L�)oeB;��ȳо�-�H��'W�xϙ���G�J)�f6zT����_� �8}�J?����n{��������ԭ7Mi��N�y��1e�Vy�ȳ�����>�侳���(�����泛|x(�Q2Z��wz�񀞩W^�4�#Jbf���u���P�Gw���B�l7j�ҡM̨x+Bo�}���"G�,)++����΁,�23����i,�	S�=��6�V�5c	eQ���ud��Q�y^1(4��XBv�(^z�^5,��L��0��d,ħF�ԉ8�/�G��΃�k�v\u���7�P�%�Y�GS��h�M<�e�Xu�*(~�<n���kr郚$z��A�Q���wA����R�	S�
��.��ĒA��Ά/� .q��C�َ�����Bw��Rѣ�oQb����shk��t�i|z�0����<d�]�ܼd���g!,�&}������{���k��)ЩP
d����q	,���ߐ^E��zi�.!8�d��m���j<nL�~Ȱ2&���&�M�K�5�A�o�U����>`�w	T���p]��C��K��m<���5���ڱ�(8p��oc~�~2:#�S���ֳ�a�5�`&�lb��}Ӹ�Ձ�0'�9�L�%���!M�:@!�ª5��+�h��.���%�f@��a����&�鵵�޸�_�_\�aFmV��h�1Zy����.�� ���!��d�]1��O�s��|�D7�;S��OB=��u}o�^�5�����)�T�%�Y�|�c	:�5L���Ta9��&��+M�;>�q�� ��������uE�d&�f��`�pGr�1Xm��)y^i̗�Ley���)�S��O}q��i?<b��o[�5���?��{�8��5��&�<����_�_�4�Oꔱ�2H�9�e��Yɜ�>�rg� ?H+���[*����+�}f͚�/����>�`Y[�WVZE�|�J�^>7⧣�)��T������J�V:�m(#��'����2-ˠ����Ӣ_)�$�X��p����G�@����(�]"N2�2b^#���� ��֠/𼪍^�/�Ns����~�%٫��!���ў���s��+q'�����k<�
f�5�ɯ���Ľ�-t��-�<mc�Ҭ
Zl�����\,Bk������,��dOD�Q�n�oxE^� �C'�j���\����/A�5���4�}��]���6�(�L%��Hxx�/~�_w/�<�F^�����!t�1h���q�>q�^ W@��%,~��q�&f��(ʬ��^(�o--U�)��v�,����#r������ҁ3���5쇝o�X�3^wZ:fw?Xb������AuXp�4�=zUCV�&;:𼥭�OH7�'�U���-M�ㆣ�r7&��A䷟��K��j�w�6��A6�2�-�*�_K������~�m�m�d4���Q�Yy�I֥R��0����|�)�v�?�ʕ=�9.�%/B����s����K nW*�#�,m����[�A�t��X�#Q�;z�E����A���^���(� غy-8ϒ |�pL!F��|��D��E�m�ߩ��e�3~ء<��_/��sf})/>��/Au�Wz���EJ�� �D�>�L��d�kh \0�g��.��V�N4zX|�[/�����,�0�9�|*��/����
޳�Ş>A�Y~�^��GHA�x�����_u�l��� �e �������1;����X�@(eB2�o-/U��"�^�쨀r-{s����]� �	! e�v�ץh9�He� �w	g�����8�������h�[ ��@��חD�j����OLͫ�:�x6Ru	.,D�5<lu	X��A9蘣��)��72��jqP�b47}W��D��~�����Z�6��ͨ�B~�)
�3ӌ~*�m򭶉��M�˚��(꡵,���ŷ�um���1�r
6">��@�h����H�~d"X=�����U�o�GUQR�"`7�2�����ӥ'��>�{�s|�ʺ~}L@�������R_�|\M�^&y��P���V��GAJׁ�m*�Cy^�s/�|�IFR)�R4���	;��;�.!��pg0�Yd����/>an����͡d�:�_�hW̓%��o�X"Sꠇ�`�a0L|�07�o����Bܬ�W�����.,I*�W?}�����2 ϩ�ʬ\�$��Q�O��x�R�)k�E�Z��ò!�D!px�K��g�K {X*�+H�K�W�������@а��� �����G������y��?�5�3D��V�<��f4�^��`�r�I@ox:�h���9wa���H׎7a��*�L������_�K�?�,̰giPw6������j�3Dx�p��S*�G���:��,H&� Oj���l�X"f����y����6��Ě�LS�gǬxbqv&��"D���JK��]��4S����/�Kϓ���/�׾\ߵ�6��5Q���}ɫ�XU����%`�Z/���_m��!8�斆��U}\C��p} ��H���o������z2��F~�]2 vtՐlX
�7�;�5m �4$��KC��I�Qa�LT�ej ���l³�lY@%)��]�
���)�7�m	��ɾ?�n3\��I��!�I������k��qS�!Y� 15
�&v��l���g������b�Q&�rh�[>�p�1GT�@��Ť_p�x^0#�ۨJ{8]ۂ)�qzy�_�&��R���B�(B)|�+��|�ݫ�������TOl�b��j"O������4���u�O���4Hf�Y��)��ƃ wfQ���ך�A������́�<���0.�|��x�Έ%�>
~����5��,��+|�a6�U%��`%0����V������F?�c��J��b K�!l���]��.��;2�n6K|���p�V�����Z�J��HϹ��L��ڛ�A�Ϳ�K�3چM}������'1��h��y��3����G�Pg	�/�+W���
cU�kQ�@��h@c)n7�	<��#����!Q���&'�Eg�1jtUH�<b����LhcK�G;t��/��Pƃ:j�Α�Go�T�2��V��5����_9V�"�+9ʨ��V{4R��p�$w�@�=��]�po�v����z����3�?p��.�󩔊Wr��D�Qmǒ�ؤ��Fv]����MF�����X��ET6Q	��h�D<jT&�j�yu^N�7�cy��_64�׵>��-¾M
���	��]�������<�5*�H3��������_ų�W^��
�A?��\�������=��4No�g.�Z�������]���'��L��/�@3?,V��v����nZqy�n�|�J��_̴�nz�`�y�r�&����x�T2\j �m>�1ϻ@-�~�PNkEyZ+E�u��3F�Uf�U%eXM^��:���_�W�/+G8���C8FTיў�h�@2h�[AR�����]Rd�+�h�!����:��h��cw`�G���Μ8�,�#͡f��h��y�{#�2�1Zu�qƂ����R2{� J�-��1�!2Z����[G_Ќ�f�W>�҂�s \]G� �{���HW~�y
凢k�PĹ�9��t[���4:��cR�E��%x�*���h���"*j�|F���uldL*�&�ڏ]�"=`s��X��N��.@��<�i ���&5�0'ڽi�Ԝ0�n2P��SgƹqT�M�W� -V5�w��X_/v\W�Җ�[q���Och& �Z���Z��EM���ژ?�cj�I�Q�Jk Ӊߌ���[�=��f�߰*��Ô�p����=�M���`�И��to��WU���������5Й�e{����;�X�U��*��c���#�۬I>K#��gag~��-/�__���[��k���g�R^~�W��.��������a�q�����p~����_���Zx�Wo7���|�vƇ��EPx]_�O{��������^C��k)#5��疻,�PV����cH��Y���:9|2�3pp��J�\�y��Hb����1��/:� �9*68Q�������Xqh�:�p(�_��?� �eç-��(�9-v�e�[e+ԝ+�+w)�ˢ�0Ԅ����=��T->4V�]MM�\}g^V-2� ���}m<Ϊ������h�%4[⎜���ݷ>�����:4��A�2��D?�f�-2A���6�b�4�	b��}����I���^�,��q�����Q�Խ�$3}�`��+����Q���w�u��׵���-�ցi�w{(u�����(ЛǕ!��J8�ނ�&��}���T�7F��ut�>V�{�1���+۰Q��eL�=����(��h�!:�j��{�a����xA���료u	>8���EW��"�b8t%yI2�u7�@C�ŋ�eD��/�rT)w4���y5�;gj�;F��ԷUt�3˓7�e5t����ɘY�Ո^¼w	�PL����R�j�Ad�L��� �B�iCs���X���='�� ���uA����0Ү��xAc�p��"����=`�Fۯ�Gős��ߓ�7v!@�)[a�k5�s2�l���W��ឈ�=@Yz�V"Y*��SMCi8�G��N!
>t
%W�gbLv&�g��~vq>�z�E�ךz��ݦ�t	�N����Y��/��?/��;7�Nސ�Oӛ�>�Q�eD��ʼ�g�ѳo� �t�0�g:��9�wG�t����A��^��D�toZ%K<�EGhb���q�2h^Leʆ�{(�0�=�]B��aH��Oa.�  �ǨЂcT�?�јDT���C'��v�{����ah�9ʏ@��Fۋy��?s��g+�e�҈�7��3����� ��m�6�����q�掳q��A3� ��ܒ�G��Y&	��3���0�ftO��|�g0L?��i��W�ܪ��^�/G1�'��a�wt4�4���ޡvF'� �x\�K����a����Et8��}:�ՔΊkT�C������^i/C�����K:G�?i����0�ޕ�nXz�+fW�O�{-֕���f��e�sI�G޾��%t�z	G��Ty��5'4�X�ǕsK��b�[n��� r\���T]��0qiyP�9;.ہ�ȉ
��3�v����
�zU�)WcSXnVk����9z=g������^������y����ļģ�L��K��w�lO��v�
G��;��M�B��&}#ޒ��}��o�2xX�����-��Y�?ld����/�=&Ա)�D�r�h�qj��ag:�9�}~$/<�G
��1�}��_v�6{_��������j ���+&U ^_��A�k��I�L��W��;Y���r��g���z͓����������Ʉ�����_sf��<���ם�%��v�Z��(���U*��M���6#��C�A>���-̵b�zE�4���n���2NX6�CE�U�а6l��9an�Lɫo��FG�Nm�c	q��O�x��n2g�j?�=������;��k�Q��Ă(U㐆�}2�RO�0�p��L�d\U[�kU�~P�WD�Ma�u��Ŗx�PǍ�d��U����o훖VQ���96 ^eX�����˺��_cz��C�W��F�d[>�]>��°^f�������iX��zMǿ��_J������@��o�r=�B��*� �|A8e/�,-�: -Ur���}�J���k4KįOc^�O_(���$�q�0̿Q�?,�|fa�2�Fqr��8+��T�x�0h�	�ޚ0E-�Efj�����9��1�<0W�E&|���붉7S��a	-��}���.{�inW�L�5�s���~��^�7Ύ��xK4���j�-|���C4ڽ���G����Ή���$C2
>��[���=Ϗ���O�)�j���[O��X���v��p@�?�����9G����b�f�<V���F�o��1�ZEb��~E����}5�õ׳���Z}�F��{VG �$�5�ry{������|�-�e�M��I��#��yќ��8Vˋ��2���п��%�u#L~-t?=x�7��Q&w�+��W��g�����(�~���@��>�@w<�4ug�ഺ2H��GnuA:w	�1;�k�/��`r0��l$ N4Ő���	<��
��W��J�5��vMtb-�Ii-v�Q@����x*��\f%���~��<��9T7>�u3X�	���(t��q�{'�2i ���mG'M�`���u��ZE��d��f�A㻿Ti��mn��oj��׾��Xl�����&qY�qC9t#���6�ZH4�$)]+z>h���q�Q=�N'N������(��mI�T�����%x_�6������1�c�.s����[k��9���}m��a�8���eg��hS��d���eE�U�Z;���t�jm>;ftqaADm� v��Ɔ�Yd�|���&^�K>���:vm��>O����j:z�Zz)/��{".�k�����Z�n�D_�q��Q��j��=R�ʈu�b�Nϫ���X"���Xw?�o^����$���FB�ܞ|�\���k_8vu��l�1Y<[�}�@bʯ:�6��f�[��*<�k��lvA���H��X�ܻ�������"���:�����ң%|���/��%�X	m��ۺۦ�r�!��o��Զ���O���y�[���S�.|z��b��Z�i�������	>V���%�};�S}���y�;^���κܯ���������5'hE٘u�-k��q<����Z�k��]G�����e��:9ץ�(��G78��R>_��B�+h�k�����s���!6#����O�\��1T��ֆ/B�����s�%\V����F�Y�/"�fb��&7@���l��d��<�U���K}:��0��ƀ������;3�AY=#��!x`%�&���i��B� ���c���u�u��zA�,�>�a��j��rqp���k���(�����
��qP��h����PslX��̷�KT��wtDl��r6��q�hV�5��_*�Q�0��.)zT��ML,�[n���K�BЇ�?�\`�g�?-l���/�Y9a��7#���n
�)�}�>�SAo4���ZOޙn�T��<' ���	��At~��ߪ5-U�<�D���ҥ�{�֔����_k��=pYڏ�s�zJ���h��ѴΡ7{8���VH �l2}������э����=����iib(��,������t���<M4������h#CV@⸟i��,����3�i=q�1E�C�P}����hI��]ss~N�I�k��Jrw"Y��Q�e�����6Z�:Lh�c�~u�hg����d�?z1G��)^����~>�S��*���g�Y�k�)�N9So���2x��V�� y}%�=IT��{?iU���Z?���B��D��UA�_nw^"f!�m2�*�2��(��V1z����#I�Gx�%D��ET��KlZp�E2��D�A�t��WgU��!���{��YJ�x�i�>�㻁
Z��<'�u��(Z'3�	{��V0��� �h���MF;�S3�鐅T���*� +���a����ݡ�Vh��2¾n\�Uc�9��$���?P�*�>��� ����U/�9��C�||!�A04��(�Q9�G��k%�$�T��6�����ɍ�����|ް"���R뒼���CP���j:D��w�n�Ի�M�X��ԛ�ݹ�R����K�)Bc�u�����!]��F�o�(?�&��*�%�k ][��R�fG:7��EK�L7����=���AK�b�����ȼ�=&Ahc/�1�:M�n�v�Hm�A����7�~W�=�����b>ʣ��'-�v��GS�cc�Kr�s��;꧎��������Q�E�w���V�zh��y_�U�j��v�"�>�Q�Y���-���K	�R{������/6p}�S��� 8���G�ƛ#�5e�{��^�����?u����u�R�/�ꏼ��?wǟ���!��fs��szM}rS�5J�N�B�7�'ST�T��
�֑�7�oy�MJ�((���-_�;��B��|p䒶h�Yr�X�]�7��#fJ섰X�F+�d��h��ae62�n!o�wД:'
ԅd(�mx��B=Ѕ�!����`�uo����}��mh�aMk0E��c��$�tl����m4���I9�9\2O:�h1s����?G;tQ���i���D��O��^��_�)dT��z�qｓ�a��0���@�>�r꫒���7z����]�����l�`�8����2�KPi���_���R�C����R��r��	�c�^V,VXcÂ{�5:dT���1��ҙV��Y����ne6�0��nS�ib�4i���A������9sb5W�Xi�����������?�fv��A����Y���m4T�a�+i��r�P���4BDV�L�:����#��b*�m9���D��b/��vO|p���0�W0�E��9,7>6����Mɭ�%Ȩ(��퍲��o�_�����Xʀϓ�kC�����2�W�p��z�fyI~j���b8?�GS�ӱ��)�,�|���QL�r�:	�8�}�հLڰY����1 >5�[�N���ߵ"�iJ?����K���������֕t�cW�~t������ӻ���$6���]/��+�vU�MVM��I�x7e�W���2a����m���7:��eJ-�x����5�d��A�4����;�JKӇ8J1Н��D'vaX�W:���Z�m�ss�U��;�Y�:(ګ\�9��}���պ1��f�?�2����9+6��֨�s'.M�S]���E�͍��e��V@��Mԣ$�t��vI�iIJa2����t���	�V�9߈�o�
\W,+z)�j�����*� ���3$D��7��嬣V���|��P���W2��=�FG��6�ɯ�^9�W�����}\(9(��0V�rQ���%��i"4�qJ̇��|��y�e�A��״��>|�E3$l<
��&��A(L�ٰ������3,�����E��\ߟ�1:��M�ݗ��zأWe��5ӭ50���+��7�.7<:(_�-�J���3�bC��/ʊ  bP�fs;Ή|]��Z���"����]�>����H&�]�)�lX��˓�o��5������R4����Ek����~dwB� ��9?�^1_��_#6��Ե�Cx��}_c����f#0S@��C�5:��拓�[��\sF��� ��;�I�����o��d}[{���J��slH{ϦO�p��'w�w�;�֓?ת�[gw��׽�_s3�ۙ?�k���1�#/�2�r�_��k��஗
!�rAi��#�k@N8��C��6aQL3<xS����y-X%D��I8� ����yn��9���ـ�p@��ë��Xkq]kc��R���k�J�nӪ��㛦7���"�<Y `�y�y���>ṱx�z�%����m?~�t2f���=�H�x���a�5qa��Fg� ���}bqK��B��
�/N���=n�~�M�]���(��\%�5�K���Zl�y"�-�̇��4��P�F#�c�0�$�*�I�ĉ��X8\%��=Ƞ��0��JqJ�CdLTo(�
)���1k�aY��o�d�[�i�9F5o�kA�?М�y��5Z��R��0�!�o�U`�/s~V��Wg���5@��i7���-�Fa_�j��::�0��낮��-|���ޥ�iK׽��<�)�+q���緯S;T���tN�M��2z�,�{ �������h^(��Q]=o[񽹣��L;_���%��wH��ꏻī��N� �z�-i�����=��qC���+��-�1�;��|��>8����y�4_ݭ���̑�j�A�1���׾�A^V����~��?����ܵ��o铽^�ʝf<�x������Q����9�#˗���E&��n�Q���kĴFw����g�evZꔈ���E(�e@�F�����g�]�֓�X�KÏ�`nv���{U&l7���&F_��!��qJաXo0C���0-M�u9[�_�-M� �pf4��V����Z�0e�qՔyɨ�f�{�9H�|$�8��c!8�f:�G�͂�`,嚤BSz�Hw�[2Q�r�uų�J"�k^W#��w�r��{���칏×38��	*��\��;�K<i}!�������&��M�c3�!�/z='}�J���Y�R�|�=�66&�m%)i�n�����:�в���M5]'�iJy��'�Y#�s��(��F�575�ܘm�,h�#�߱8�n�ne������,�|�e�S�%5�λ��鴲vޙVl���8Ӣ���]�Ó,���FG�P�*����G��>ߘ�@�{�h��3��C�ԉ-�}K+��(_���=���Fӣ1Ia��Q>N��r���d�V��{���t�ӺE��w�Q�u�l��8Q��X�3����U~��_���e�9�X��u>͐��1�?j�:�f+~Y�|*�o�,C߯u������M�A�������c�|=
_�,o��W��;�D�Y|9��_���KV�i�vz�V2�1Z�ܲahG}��v�<]o��	���_��:��؍��y�
+:�<Н˳p-�ǥ0w��%��X��h���J�h��;ȗ�A���,?�����@��*���&��)�f:7�ea�ސ/�^_Zj����C7z2*�F��/�^:�;�D���㎙�Ub �
l�W��2Hnh�Z4b��E\�@��Nj�L�&;.�L�p�3�x�q����.��!$��%��W�E��[��>��C��?�)r��!��/��ꭚ���v�YDo4
���&��	�v��Ѵ���]b�He8��M��7}<���h,a���$�xl=I��QjT��<�э�Qh��j��Թe��X���h����ɝ�hc�F�^�xΔ^�H�:�8�2�w��Ι�_<hR-AӮ�fn�&̉5c�E��R��(��G���B�z©\����]��F#Eo8ANb	��7�^�8�)������k>��l�㋃�FDY,�$��>��-�r��[Z'���M J/D|����!=f+�GW�R�K��}�~�#�%����� ��R}�4u�])U/0�j�lq_��7������z_�ˇ��ʬ�R�N���R�u����w��
�^��e�/�`��.7�<���J����7�D)V�� ˄�-Q~^`���v�rf.�Ҙ����
W��	��P��Of� ���1�;T��j�ޥG���������N!��|�����`����M�̯Z���=#������;z�͠�@���e�U�~��:���n������1�Y&_���r]�w�szt�����~�����:�ETԻ�����Pl �?V�u���X������Ɇ��l�y�`��/�_N�ٰ�hTg�&j��y�����k�����"K�A���9I���Ĵyô��!:�.�
Z�U��D3�9b	����
�b^��m_����j{�p�F�͒��uܼ��yu��=�Gz&��K��Yq�}��3Ĩp�U�3�e��{����<�DE���P֟��BLn�AT5��Q��U�Y��.�L6�(�K}ٞ�ӊ>���-��9�����/׿���d>p�-���.%����_��$agG�R����~m��ae=N9�p��N�[N�#��_����C��|��s1?F7������{�IT;p�����KD
������PPx�)׈<-un��<~o�	R�C&u�ǉ��ރ�O������x�3�Q�����#�2X󫢂�%���5�W�q_� L�:��hic�zC�El�����p�x�2���Y�W����*T�H�b�ؤ���p��Sӯ ��6s�z��D�<EO����$�Lr��=�^�BO\)~�Q^�^�9����v|��oq��}�~H\�b:E^�d�	*���|��j!��q��Z@�X�ðb���dXXP3�n}��rf�
+ZL<&&}���ctPq/\pV����|�POƙ����H�||!�"f�3Ɵ��P���F����C�]w,��@Nݝ������W�����=Jy:$������F��jLr�����kH�D^9������:�o�kъ|w��nuk�듏�]q�.�?�T1���w�3�඙d�����"{����i�2�6�ɽIŊ��WT�J��|4�'vw���?:cc�>1m�ڳ�������9/���ݵ����2�c��4|o��r�������~9_#�����L�˂N���>����}Y���Cg�kW�ߕ��2o�u��k�Z~M��{�_�'�����e4��̜�O�����gi��s#U��0��@�M����yڭîZ���"�����[:r�(i}�KF?���HF��׎�v�?ց�*:���Ձ�#�?Z���_}��g<��wȠm�O�Е�} ��
���m��Zkd,�@�b+̯r�~yS��Y�yچT}]�֞��&E�s��r�WP�����`;R�R{��
�Hg�3)}���v�r�!^)� ��;W�wt��,������W@���VEP�X=�71����h��-�<�
v�Ѹ�Pq��&��+��4�8���M��Yʥ�jiI=w���,�&n�rfU>�Gr�c,e�n5e7�+_č`�����[M�k��=L��M��ʇx�kZ�3�~�aҰ��\#��L��I~��5���)�(X*z�=��ܓ���q(������00�b�k���C���1W�
{T��F V�4,:��͌��|�V�����4�G��5�W?�-<�T�(��/t���IB��K�c�}"�����ѯ��b_U_%�ך��m��;��k��\+N��^�������|���Jed���E_��^��q�[��3��f����-a�Ll��>�<�:�6��<zp�*�b�]��+�+yʍVO,��}ix���r�R�"���!�H�
v/�!�8x$�?|(G�K�W_cW�o��m�������*0�����Kx�ľ��z/�C��!YT|���N�Xb�4��i�ԤE����D�<0����B�^H��s^���=n��/UU&�����
�ա�� ۵����^��ql	6�O��l�5��^���P�Fɣ@���y�h��5&��p��-_D_���1Ц��Nr�pN��x�����Vr�=N�����7�$ԩb5^1��&�0](ע:�����V#�׵� �cy��藮�����B<��̿-ʱ��֍���〽�(K��M�T�3rs1�YL}�6jy��s�ѴT!_ED.K�a&K�&z�+��E��M{�"�%5� kQ��1�Z��0�?�^�0Z�U�~��wm�x�����1�h��c*X�b�%syޡ��n{_���	y�|�ϩ����T��L�j;O���ſ����~�O�k�i|����%�SG��_�rUq!U���m���Nc
x��Q��G���u�U+����-v?(N���@�B�)V`Kz�::s.�n�J�%��{�pJؚZ�G�%!�l��ͽ�pT���*�:��պ-�������Y��~ۋ�m�A�9ı�����s!�0��>��e2D(��*���*b�kL I� ��ZH���h�~S����U����˹� x2hy��;�Uð>y��{�tygӽ����I�{�/��|Q��_��ީe8�,X9�j�h�L*�B����쪦�6Bm�0þkS�G/SI�KM�H'vh�=G���c���'�|6�s*�\`/u�ҥ� >o@��&*3�?�d��G��t95��$W�h*|&Yg���=�9��$vhc#�x�W5�Eٱ�}~��,U�ei�[_���wY����r�S?[�'�1���'y���:3Y���Wm��Dy%c�}g[����Wߐ
ӁJc�ӂ�N��h�d���.�yr�=�3È%Lr�%��2r���F�"�A-��娞��'��2�st���'���
R�m�d�<L�/)��}jq��2z��G׊ib��z�n��;n�q>�{�N3R&������%[7S]�u��jZд;C�K����/�CI]-�c4��v���R�?Z,Q��H�= �Ώ�������9�o��ZV��ù-w�~���ESa����p6z�n.S7����»Yx_�9-�1B�0�\�db���*�GaN;*����[��z�±���h
Q���č`�Ǆ�B,����8y��p"��טN���q޹e^�b)�����s6H���|�N��~՚������m:rYp�q7ś��h��7�8q+A��0x�{�J��:g�	p~=� 5:�=��o|`ס�����<��B�>KBO�&HKW�=�.�Di�R�X�~���R�?�N�g��]���p
���ܯS5�m��Gh�Yy�>���L�Η��$odl������x�R_��K��#��t�Rk���ɚ��su�^��<�\����»O�������ѳ!6�l���>&�������?t�|H���"F��&ד��E��q��n^��=���כ��_�t]]h�đ�&�����3��3ܟ�Iie�y�}��RՉ�3J�X'YOU�m,���Z`�*h��8[T���1���0n�7�:��`��p���^�&��D\]�q~��:x�Y�ȸNj�e��|����\)?��0<V��l\��(��#����:I�!�r�w��h�P5l����*��n<�xjF3�A��p�q�S�M������r"���I�釾(����q���O��r���2/���kǖcX!�ypy�����U�W����jTX�ӥ�s�;��@Y�H�?�:p���b^א��f����JV��@ja��;��{��Bn�/h ]�d�Eay�z��oY:����[��+E9��h$��w�[���G�ʅl]��}ܽ��mz�sa����ֶϛ�ef�
��#�/H�a�UH����n�_���F�U��#�T|�\�����V2w䋞�W4�\�ϒ����w>�ٚ�j�\j<K!�#�@���XB��ho�]�ڻ���a^��C��
�N�V6t�r�Y\^���2�a������B�V-P�l�	S��������5�P�s�ic&�.W��(����t�P�+�E��P��!Hmf��ߌ%^5��D�o]Y�}�r�� ��$�ۘ�"t�${4�����E]+�f��ƑS�r��pp����~�Qx��_{�|�����ЯT�ٱtE�	����;����➷�P}
�Z��&���Y�]0;tԨX�3�/� W��s��=?0k m[�쬉oc�>���(���P�=�x��Ȓ��]��^�,��c	�t'��
,sk�螕Rwb�vy)H'�Շl���昡Z�y�y-FY�Ұq5�y^�h.'�ҹ��i�κ`2��Gay�n޵n���t�(�Uk}�/���u�5������v�w����?�l�m;��Y��k��wz�5s��V���/���pΕl�)��P,�R�rJ�nKQ�!W���#��ȃRq4����I�E-�5.ciR�0�2H
�6���&fSe��~w°K<��L�Rũ�"���ޤ,-( ��ɘ�9�ֳ\� �*򫃂�.��۩�� P�䋌tV-]�����(d�7�ud���L���\���v�V{�T�+�^	���A�T����/���ף�o+�A������#H��{:�MoS�T�⡹��4G����DU��T��(�`����Ʀ��r�<���|V�]�ec~UY��4�.�KG�a�����?��lX&�������\�&����!�B&ÊgO����u]��%�+�
t-]&Xk+�1Y歬<�%H���K�	P��B�Sܪc������=��|3�14>��F�kw��<�����]�}I��G��Q���|Z���*��1/*��ȟ��z�hB:��g<���~�_kB�_߻6*�c�/��J�e�>��׶�A�����u���ԑV�[�}���ֱZ��]J������?����|7�	6�$?jr.�C�˄�ݏ)��='M�%�Z��ӾV�t����u����ʯ�AT�����&��Ny�(|45�u�.1����h��R��9B�̦b�P_�����(/��T�����`ʈ�˵%��O~�˵��i1�y�m�\6/�|�D��0�r��T{�w���A�a,198��P%�8��ͤ��!�{�Y�V���z:���R,�>4�Ӕ��%���9s��q���V���&��H��櫟�\NM6�B�EH�}/-<W��d��em�*�Wx�2}�'���� N\s�p݈6�W�k�}_��ڢ����}+ZY��f�Z�ځU��<�<u�ϰ�x��魴�{���i�q���|�&GQ��\Z9����Hy� �(�4��Y�p�X�<���L�2�9��/�s�Uc}ɧ_6�M�w��|Q���{����ʹ@��
�VNI����3�;����*�>F�#���E՘���� ���q\*��s�_F �=(��e�^�b1%>�@��CͻHF)C�f}֪��?��j͈w�(m�pG��7ƃ� <�N�X�D�~T���&Z���!�*���M�Ԗ��@��p�l���BQ���u�d���?�*��7D/���s�y��Rn,���̹��t$�R"�
mV���*�h�����s�F5�����t,�c��JU�}qb58��.�+��c������W�=�{ ��?+�.W&F͋�F��ڲ�T�Q.@n�K~�p�Y"#f*ҝ�$��+����qwiwm"Й���CQ�B8�_�ʘܳu'�y��n��\;,��5�
^Ӭ�E���LZ֑H�����4m�?��u��{�%5�k后�C%�6�H�i�6���_��悽(ڠB�E���t8{c@{�+�H[�Ɓ	@�Z�}OCt)��>S�.����XH"����$�缅�:�Ë������Mܻ!~E����c������-��*>�O�]�!�YZ9 �TL��]7V�
��W� �6�@Q.3����
��巗5��O�r�0U��4����U�Ϫ�-��R�B�X"r��Ru��<?��z���
ɮW��Ҳ0v� =���m(��h�q��k�\� [ ��A@�g���5��1r�.��̡ޑr���أU�����k�jw��e3v�������7]',��Y-uc�.���ѿ��..�1hU�C��O��x��qs�����wdOu�����3X�Q��x ��X7O���u��y	��# ��w_� °Br��X�����7�� ��5>㠵�������_Nt���5��)Ď3�"<�[pv��n�	�_�\
�6����`���>iq`��l��t�>��	��f�q�@qj˼}��Q�c���hZ��2c{~�q�qջ�N0޵�Z}T}�%��u��x n� �|�_�
/�e�Wc�W}�i?�Z}���s!�y[f|��?�v�J.QG��r�%(~�9��B�����B��8�[�楶�tåO���I[X�!$��
�bƽ�k��b�J�,Fq�Lw�ؠ��8��4D޸�ܜvH |��q�^繼V��Q\B�F`��V�M���S>P��]�E��CHD;Vxq�J���K��^я��9��0��ixlHpdEn� �(�p�-��G��y�_�x��,k>&�.q�\����K�C�1�UsY�`�pE�A��׌<	R!E��<���*�MV�����wӪ�y��9b��P�@�Kg������͐���O�sw$�[�ԍٓ5��F�Ve?�P(��S?���b@��x�`����lg�
��Bz��_UӯJjS��W��A�ۦ9
OݙYX�ʫe�T/y�\k�U���K�l�1�u:���+�E���9o�֧VA��~�N3TWk���u,��h�C�ڡg@ϖ�VθX�0��������D퐹���k_�0�nk�Rc�G��I=H|���r�&�Y`��H�v����6��ͧW[�����MYu�������0�}���'�}����:Q�4K��6&�L��BR�ע:Z�S/$�+�u�� �Ɔ!7��5��#��+�q�;�G�?�!q\jJ��*�ZY0��y���%Ը��,��M9̕�:�Y1\���8g&�y"�-m~C��0U���y&~��y�K�}i�|[�\�铲� �l['S&vk��wk�\n���EHi�M��'�⬳:�s�lOK�I4�V���I�/��
�h�pߟ�Ӊ��Wa�?�Պ��4���eJ�%�N�B�4B8�9�g0j8_q$_e� _yE-_����TD� �`[�޴�\�w�>%_k��6J�O��.��Z�����*֞�I+z�>r�Wta9?�f�И�^�s'�����*T�z��a)W\��&쬲{��B�r�X�:�S�3S�����%���)�Ⱦ�7?0-�ѨQfR?���%]0�E��*�M��г�ϭ��	@�@(�4�˨%��z�L|��D�Nnj!�;�!�5���xŧF\>(����r����oR�L5�n� ��Z��>.(���vܤ�\S��-�1��.�āq�q̇��a�=�al�~�&�	1��@�s���]�=q��r��`p=e��V%(�&�EBC�X���K�r�BdMf�����ٕ�K]˵H�`�[Y����	�z/,&�.Ƞ79�q�"�=�s�-�:j�3h�υ;�|������Q|Y�UB�@Q����z���x����L#��+)���E��v#�L�l�3KV��]�׫�� ]�'�!A�2����^;}�k�[��档��ϒ�kW���#3��@K��w%KjCدN/ѐQ]�jA�w#�ru�G�������]�L�����f�,��Ӷ;tg	�B��-0�(T ��4�b�D���b �=8=.&O7�$mP��eQ���v�,{�Z���w!��,ь�/:侈��%���$�x68ǐ��)�pr�68��F�0��.�?�No׉$�̓�~`d��,�dq��?F�J-YTcL6�8�����\#G2m�3+����feL>�e$z�0�D���kɉ�*�= �U�M>\�x�U)�}m��D�<ԥ�sK{�FsI�*��ڻǃ�<c�M�E���pA��D�(��($(�C.��%�]PF-II8p �7*Nli�&�3�M�ރ��T����鳄o��)U���`��c�e�d��T��9o����ه��.ie��x�r�u����)���t��YJVԑǠ�%~$�y,{_6��=�__�͏ʁ(�����1�yȊ��/&-LI�#�)r�'�_ՙ�\oM^��ULl�b	v�j�d��I~y����je�\;�k8�F��P�@�i��huAk���pt�'x��DS/�tm��Y�aL6چ�e�Ꮎ��ߠ_�jZ��)V�ɍiW1ч��Idf��]��(�4�w�(itF�h _0گ�CQ�a���{dN�>&j@li�~6���"�,�ی(�a?|P�Bݦ@/�6�`r���r�/>.�ׅF�8qǺ��V�vN���C�-[�߈�]���Fޙ���t�k��g;��(ɨ��w�6��֘��d����L�s`
�.���d����B˽������ܜ[U��;=
�c��w�)�r���KG(~��3�������7q�$x�Z,G˖Z��	�_k?T����{���h����y�?��O�������<٬�$-G%Ν��@��y`zp֍v�(814O�N��cre�#%n�E�L�1|�����;L���װ�S�Ao����� D�Wt�h���^qw��fr�2�q-�����2�60�C�A\f��B���\����BPw%]�t7$�W�u��˽����Uo�tn�r���rQ��|����Y�D���ה%�fU�1Y�`�*@�<��6^�c#����+/ȅ3N ��ԉ���ZYᇽ�]�����U�Y�k�,y�uc��g�7��T,8oQ�Κ�{��oT�,(�y�j�����Dx��uu�hJo��e�٤�����q[��k/��s��$�l�[�V�/o��������%��s��������P�\�����4�e�r_�#����8_ń���حֺؙ�8�����S:���x��u���s7l����c�r��Iܱ���S�ն5�=$�7g��e�y҃`��㪊3A,�B&$��0��)@ט���>@��I�/Bfյh�!���^�h23��Y������|&��8Б���w��\h�KD�-(lw	�:��� ��.���2�ؗ�M�&��>>i�M�yj>��k��\7�-�~�)L9����X7F*/񤭂�zi���ug�y	�>��|�^T�p�֙|k�~=X*�D�d�\��2�Ң�������%�6;Ӷ�;_L�ϒ!g�Չ�>WAf�ޤ���K���}}.آP���  �.j�1P���ˏ�����]T.~Mt����&}���}��_������%���m���y[{2F�jNE�5��8�|A�9�5N����q�L*߭���:�=5?�%~D*E���60���ڥ�:>�e�0Y	�e�7��J��.�%�6k��6:������U���R��Av.�=ȱYAgO����ͫ}��i�@���f��0[�Z�1bjoʦq���|�[�ÉE�A[|�.��Y���(;���r�s�Y�]��<�	$4pn������^�)��C�ۡ�h�R��gi�\N�;�K������ĤPK�����[Z>�J�8�k݋)�_�I3+�w|jޫAc�q�`��/*X�~`�7'Z�X"bb�Ԛ�sb�q�֨�1��C�yZ�b�j�(|��
����n>W����.�פ�Y���Hŧw���'��}�N�<��o~ĸ{!�%�u7½���c���2Q����)}:����o8c�Y�9N.������i'�ZĒ&b���]|Y�Y�֗��5P^��G,�{q_��σ�V��H�A��8��l�Q:|���aeh�OG0g�%�V�t�ɵ���c7��̒��Ht8��|��������j��x�5�̰�e�v�#X��6�YXe��E����`�]i�7�7/5�+�z�ڑ������X��Y]���"��.�u�qp®Gw�C-~A��
o�K�)\�65F[ZY<?�:����ȱK�ω�q�R�^��N�n���}B�n��4}H�]�8�F��W=�����Ou��WA,rٲP�}g'/k����0~S�mBR�WTT��>h�����{z���;Jlqԉ�>�#��*��6��5�{�
�i�Z��ݠ=�# �L>p�nC\�λ#˺q�(7�0�mH�Ƥ5�\�^&����&���t纋#�8y��SG���V�D��&���^2����eQ!۫���7[�O*���)��E��@����+rj&p)1)U�{��5����L�� N;-���>q3��gՊR�6fwl��G[q��Ea����<��K���Z@*q' 8nk�����޾&�%䯭��3�u;��D��z�6!�Dַ��n�yo�y �4�^�B|��ȩ|�]�Wo8�{V?�{7�G��穩V��y,�e�:��?��<�\��i�C��,n��ͨ{�Յi~��oz�ͩMن��I�:l0�T�eFƵ�#B�g���|��P�59o�F�`b���!xb?��?�?����v��Va�7�O�+]�B�d\�y��]�C�/��Ǝ�Pj��7�U_�J��1��
�{��H�©p��D�ب��fu�k�.y���k^�%P\�m�����o�;�V})�_5R�z�ߵ�Cy~�R�r�_�_k����n��=|�n߮�}e]�*������<+OƗJ˳ڱ3�n�L�[���)�2�XB���D�K�0����Y�Ք�H�&�J�!��ڵD��M~Ox��c?�>c)�=�c(
Y�=tf��7s%xw(�`����~ɨ۔����I{ �������4q6�Ⱥ�^���Ψ�C������6,Qم�yYc�?0r;�+؃���?4a����:L-�`��[!اi��uD4g����1����ܠ�����"�b�G5���G[lml��������X(зw��]C̭���Zm�+v_����[�X�*:�K��;kk�^^�km{@e_��!�%�~]�+�����N3l�N���W��!�gQ?��4�g��m���[`�S����N�g�n� ��'�e�|k] �ƽeÔ�v�a�u�� E�Z%<�J�^5�3J�|�N�Z>uu��{M&�;�������������a��  �Ӳ#^���א�aa�c��t�-~Z^Ű1�]�@l⽐�E0&Td&�-�d��߂Rb�$�1_}&��� � �\:u>�ˣ��G A��(���c1v˰�>x9>L� ���a4SIΪcy`��9���Z��5����k���zp�8�U�t�J lT���������y~�i����ӎy������ql����o�c���y�������̅w����=/|���p��'=+F�;�'S�+�s_��G��=+����Z~~䬞[����]j^AH�@[*�bQ�2@)�b��5B�܎Y0����%��mwxE�2�LĹ�_�!����,���+�g��[���AiG�B����	YoG^�<W|�[4��@�0��ܭ`rs�V�
��ǵV�u���u0��".G?�e����>|��;����fӰ��)�F6��R��\R^$Jp.�_�jp9:,�4d�r����z�5;��S��J���M�ռ�-�����ru��n��c���Qd0]Z�z�烰K��4�}nl�����i{���<f���V��討� �X	h��(�VK����ߵ��Kř������k�d����לc,�c	+�Ƀ�D�s%߹:�1nh7��f�q��਍8��g�B]{�1L;�7$��]�G>����-�^�W�� �Ŗ�����˓�a��TLՓ�L�GI��%k�[y�->Lތ�:�4_}䧸i��_��G��#7X�.8@)$�EنA3$Xc�⌰L�V�� COw�����D�#��@��D����
��i*��@jf.�/�J+S�dż��tr�$�}8_z���7L뻜���`���5�iv��7`��@�r��Z��4�p����]uTi"�h#����;9b^e���1�U�D��,z�Y�훕��Թcv84q�r��u�B(&��Q�<=9r���9ǯ��`�ڹN��j���p�3��q���ɥC��7Ί�t�KM�K��l���Y�	S���5C�a��\���%�����v�e���a��J,� �b\�-�b�3&����3�׹�Q��1��l��/���<BN|5&VGow���c�t=�)�q���~������[�����|ۚsX�\y�G?�I�[��6��Q����uȒ�J��6w�Ҹ�)�FqrRt�2	6��jh�[L`�)��"�����ɃPπ�kBE{P��=u�NmEF�K#%��Y2Ӯ-�Q<�ǥm\�b� �9p�zA��;L��I��G,���N�bI���DqbF�u��]QTL�	a|O0:Z�oLK�;���!�bT�����_(��fk�2�&��YM�i�v'�1
��ݯ�P.V&����vje��z���D�t�u��\��	�^Qx!�5���]�eX%�K�X������2F������O3��>3�"\Q�&NU��^ LAsO<�T ��N�{X-����������i��ܕ�h��)=?���S���9JNu���Rj�p����7�<�L,yFNu]o��Ig���R���.z�=��-W�]~���l��%~[&A�	�9���O�!r�k~��<����nN�z�V7��ςR�P+�j�AK�5T?���͵N��uR#�#tw&`�����m2���S�'�A,��v�/P�����@R�eG#��wn�k�F�w)�ռ��ib����;�^���n>ˋ.3fx��}ԕϹѐ�sǠ�7�5'T�c�J��$��>�5]�i��.�6�6�Ӹ����\�Q���zx�ŉ��/�Wq�	�U|��)���;�a��=�M�`���͸�C�{����vmXv�6����s�B��j+��z.������|4�
��]��W]��ϑq��x���i�������~�D)O6N)'si�KD�0g���9�K�ɨ'��S:y�XY"�L���TK�P�k�!��P�,���!�j]��E�E&��A�Ҋ��2Za]<�I���jh;O�Mh.�W�W�aC�����Co'qK��/�̅�SW	�)�/�qu��[�*0%�J1y+���D�3�������c� z+���U���8[�Ҟ�S�n���ΙvUB�5���t��[�fx~��)����Byws�9~�f4 �8�3V��,Vˠ�ڝ��4��\u�Ri�K�U�J�R�h��y�f�p3�ѶS׽x`�,4�&�|��h�T��30g��VO�qJ���e�q8�Kt~�S2�kX����s������=>�N�3��I-G)�'S-����g��z��U�Bd�l,�����O�����Q�U���u�*������ӓ��8<�H��	�>�`,k��8Q����&���ì�x��?h�n׫gx��j��4�x���x�H��"n�0���K��c�Qz,8�c��!��>/=Rz�Y��P�K��l|�� u*U��l�X�9��͝�/�cꁄwGw�,����kl/��VηX��PA+�����^S骾	���_�q�"������u7��hб��Fрv0Ō��za���x�bvq�s=wx�Y6�3���|u|_�FM�:կn�k ��闼�;��3{��.������qj�Q�s�Z��h�Y�2J6H�3W���xr�b����Q�ݢZ���.�]��Pq�,��������C~Ԫ'7�����4�W�</��Y��9�cG] ;`#گ^�V�[=�$.��y�ً���c�wq��?.\������PTT�߻�v��F�t������ � �hR,��]�~�zC���*�[y?����(t��)�d�\���6yL{��ὦh{�}�U39lL\�!Xp�f��um�)C�0�_��$υ���a$������J���z�5�y��C �������n!�p|p`��oF�Qp�L�u�����Á�hx��{ +�~D���n�xaP��������ai�?����;�?���E�Z~��e��%)0'���8X)��6���,��ڤ�Vޮ�J�\����W���A|��^���CfA��w��+��,�O}c�r�\�t��2Hp,��]��|]����c^�<c	}��f-U5k����~�\�,,�.��AEg����ms�iN^Z�3��Π<�n헙 �҉j����W�]�eXA4D�}�U�	2ާHK4������=W��~��ǃ��T@<��q+���ʺa�Эoz�c}9Py��9�jO.�6WABdR�'~<��ey�F��1��f9p$+��t�)9�F~�6�	�༞ʝn@M~�:Z�3؉3*�.���IU,��84�0r��'��m�� �m-����\�t�	��đ���+H����:�/��f�Q���M6$���eJ�+�t`#�;�2��\�[64����4_��?2����l\����!�\��U�������O*;���#Y��������g����{��xZ�6]����Ԓkj�>�n���s�QWp��1��n��>� ���|��+�t�^4��&ku�]�5S�� ����E�wg+8_"�<o:=�<���J�zt8X�= H��R8;��u�0��݇�^D����.��Q2�7r#h0��"J F7������	��?�(fsl�f�hҜ�ܾN��=Xv���� �~��sR�Ju�����tl�Zf�01I\���~3R�V���g���uǷ����yl.�G/�3Ad/ �	V�u����Q��{5
J�&��E��(�ך��h��ߺ�]���_�"﹚N�:�k��ͧ�"���@�{rV*v,��K�q�c�	P	�W��_e�E}��k�ͨSJ�u�IKkї/�c�i�%�D����ݵM�=~$��!�3�����u,񇚶t}����b�����)�<�$F����F ����"�8�� ����b���V�����m.M��EW?�� -�	��������&J�rQ�3�/X�_{�>���׈���r��yY��$���$�>b\O�0p6�z������}�<�k:+��e���;�_V��cq�uC�OR�����2)�>���Y�7b;��/�zb���\��a[��G�M���H+-�%�N�ڳj`��&Ml�s8�e��p�:�+2sJa׾�Y|�8s�&������ct�������2������4�湯m+��UQW �u�&�u�3�h^��]��?�VR�=C^qmiQ� �cDu�s��1�l߶(sq��nmڕO���8M� 1�����y\�4� 6���Q�s|7�,�q�]2X�&�V<D����0Zmlh�w7�$����v��!�0Qnȁ����I?H��ÔjN�ٰ����H�4�4yx56nPT�|�-���$�f-r�Yy[B��h2�Ut[c�5-�|\T�+�?��,��;�q}�Ш\?�|�?��x�8���s��B�t���C��^o��W��aU��.���������{|
���K���s��=�e�1{}���C1c�O��ho>�GV�m���Ԁ(�R13_w�W
������<���Nɛxi;��e��YV����nfz���!c��*Ro��.A���ڭ.:��u4ݣ�T�ko�g��5qrԒ��Bl�U)ή|��*���(/������KY���m��M�<��~R, <��Їw�Nz��sծp�܈Z"/[о)��/�ҝ�S��JH�hs�A�0ж��\p��9�1S:�M��Kq��D?~���d�h�\uC��Ð^u��S�����^�b������x�Av�0o��Pe|>�U����1[�G<uȷ����D����U���#�B.�9/��+�rp8��`��o?�]������诋�ǋ'��6eV�;S�5(j�K#l7���]�Z~U���,���8�+:�������p��nm�>q���G�Lm��s��5�v�G�SUu^��|&r��X�V�����ǪYN%��}�0?��D00��6�h�A��P12�<pI��U�-�s�j��q2�X30��Ǎ�mh�4*9���z��
@wǕ �%��`�����}>r���Y):f�H6(*�ӷ3P�Թ�����ה��8#�A߻�j׷�o�����:oo=�,�v1wZ_��r��{9X�[n��O̸�q�Q;_��;2O�ǐ͘ʞ�	1�3�^�fǴ�sȱ9_��WD��̵�p�[����)��E��_F~o<�_8�{��7��įOj�7��q�lā���s�1������;�@:�CM~��ap��}6uɭw<�6���ak�C��` v�8bP3^-B/�L#�QxF�$h�1�(�3F��V��al'	8e��Ƴ�"����Ή��z�x/�]��7�V=| ���V�x�E��O�S%�d�/nK߸�%HJ�������~]��0v�\Qϓ�H�?����$]g�ˉ��u޹�s�g�[S_#�w하�6����/���>�^���
���|�货�N�w�
Q�?\�C;�o��~� ��y��d��*
���7eT�0~��*k�r�Ҟ_xL��uB��L��i�GLp����y-Q�R��	��-v�8�p}�J��F���m,nI}��dn#�+�0sa�����C%oŹmT��Q��N;I����<�E��PB�VhQZw��#~lBf;��9�ݟ����ai>��<�{�SV����.��j�@�N����u�Í{<��7E�0�R{C���/?Q�B�-=�W�ôN��@w��L^��%L�L�>�t����Զ���N��B����u�����
�����9_����S����C-�@kY�rq����w��1�B|B6�B��ݠ2y�@����k�ω����~א"�Ɣ?�ԯӼ��,�Vx/�aF��[�}(-��[n�&�fmJ���� ��w��.���[������Q��-<\-�I��� b�zZx8��� \�ƳȲ����>c��,A5ycO�:����q��>;7�|�a�
�ժ�L�.�u`�w^�)h��v ���j�ȱW1����嚐fE����!�G�.@�(�8��R�LS���8�2�|�޾%s��獽$�!?7��&N���4po*�$u4���_0I��~z Lׂ4���ѝ�Ь�b�Gj�"�>�<Yu�\3�!J�nf&�ЖA�z����/L�O�J��i8�޾�XK�d���I~�t` %w	j�	���t�Z�u�=���7��{�Fs}-/�~�(�m����(
�(�ng���!3J�M�Q�q��))�A�h����6ctƀG�JN�I���
�*��Qv`�y�}c�i\!wa^�Y*�|�̊�kt�8j��agcɸ�y����[�cy��G��pU�$��}x��y	����_P���gW"r�0�ڊ�(z�|쉐}/����7�&-uӼ%��H+`ѯ�����9���d�e	L�<��n�rB;E���#̟����q�2�p��eZ����
���l��Uy	B��K���#����0;`b۴�i���ŷ��&�-N��(�c� �通����K�L�Β>@��Dat3Dp�CgInF�3v�by%�ii3݈�?�U����d~U�me�4e���9@�8׃T4����y��T� �Y�2��H�NkD���3�4��,vl6�GsG����ҧcoЂ��a^�%ѥv�R�K9�9��l)��. ʌͨ�/w��|�3��H�����Kgx�����5c�e��/���� ���������J�_Û��.P��������ޔ���7��eݥ���9DǾ�_�4�k���$VG�� �D�Ԫm�	�m4���ا-�V��c���[����Qj&�\>MZ~�z��#��6	��T�(�1I�+�GA�4�n��)�DPxcz��ѳ����`|i{0�����w��;�Nr��@��8g�D�+�s��A�}���n�թ�N���>��iA|��4�a+Ď�&�P�󎗯^:g@;
�F�@3^��1�,�jd��I���|r߱Ȗ����[99��p��F�H1�$�|�ԯ�����s|��4*�>����ރ]H{��yK���3���X�p�0�En��7�!y�����9��0]�>���2/�XwI��>o�-����Ȫ3�p����ݽ2���e�i:�m�h������K���CwJ�iH�4�cN|3�J1A[��f�U:��Y8`V��:��FC#���.��w-ƙ�Q�(�w��{b���?*�4�UTT����k�#�S7]0�j ��M	p6��k��z�?����wmhuR����>Li�6�����;��;�^J��!$����>4�|z�R`���c������[�^1�LS����}��pM�ϓ7�{��O�DEot�?�L�?�zͺ�K�C��x�,m��ĸ�6��9.�$���6��M�F��H�c�
�����$L�Ƶt�K?�:t��tn��0�.e�6�����C>;�����Nz�f��N�3��Hf�V|y	���X{u\u�@�uA,E?�ȼ/��9y�z�?��^���4�-���ْ����>�1yx�Z��%�nQ�V���_5��=���h��&���}�>���V�]{��_����ρ�S���~?;̟ou>���;����d���
�4�>�(�i9���ϫ!U(�I�=o�n�rx�/�y�
� ������å�^��m��K0�������&��h�Ρ1)8��
m��(�Mfo�ۯ�fơ�c���wN�aȣ$�8�m��Ҍ���j�����0������(�]��h���8mƕB׆2M��J.l�x87��ա�]��:G�g�ZX�D���j�ʈ�������*~xV�0��tH}�Ħ�v(�q��G>�o��	�l�h�hР�u(>g�o=s�3���X眃��9P8�y�_��J��,c�н�f��m�-�5��[����My!��*w��&��d~�zr$ԑ��,S(y˨Z:A���H
a��x9��t�J�sX�ܯ8�^l��B\Q��U6�h��+�.�~	�đ���������Wh�כ�ӄ��a�1��~~����Lo��q�C��l�g���-� �#�"�t�}���Gth|��ol�f��������QO�Ѐ��b����Wx8�h���H�J���_ދ�������ݸ�7+�ǝm��<Av��*��)�x��OTG�&��`������m��������d��{��7��k��3��l&�]��
�c�g�����������*k?Z��#E���`5��U���+�%�k��5wW�r��9���y�u�O"��kG�S���8�s����ʼ�!ڮЃXBU��yJ,��ꣴq���S�& s����H����C��h313����VR�l���ʯj���w�Y�j�V
��52>}!��t��/��I�k�2�m�ڿ���\>����2�i����ք|O��}������(�����a2�w��"����`��0��1���Z���̞���@�B�M�A�b�Z|\H�bߩ~�u��K������s���D�\�?�V׊ cH�|�V�"К�i��T8�P�+�^ճ4��h��#�m��3�S�~M&�v'����'S>;����|`uM�fk@A�x�92�	�bBҢ���-u��;-8��.<Aׂ�����g�,?���z�s0*Cر�}ۄ�m����n��'yp�N'��)�;+�n����=<�^�*�N���9��|�~i���p_V9�1����{���	}���VF���1[�>����T"jd8[%�q0�>��M����e*R���ݞnk�e��W��y�p�u��U��ܚ2��*J���x���a�Dy
8S�]-�e��E}�u���:K���y�*}���5`��nӃ��9�#��H���?��jq���JC3�蒮�%�.f3n�����:���nA5�({�,��8p��*�H��"�a쭮؂�w�8��X�w� |
ց��7e���;�𪆣�q��.���߱���!�.d�g�"q� z�1ѽ|�?'������m����2�S��uݹ�hOV!^�k^!�rg#���ʚ?����K���s���'�F����A� ������q��Mk1����Lt D�P��=5uЙ�G��e)>��P��Қ���7&�a�?��X�-d m���fa��l�+ˉ��Iwۗ����"z':��m�%�WU"��x���憆����9=(��:#k��kd�/b r_�:� �2ɫ�����|�lKNw	NO��"E3��9`�ř�#:��� �Z���$�n�]�;�,c��V��Ɏ�"��n�{@'��Ʊ[g }o�/q�p�5��3_,���1�X����������^i���v�t��|L<����}��'w����4?��y$r����1G�(E9\i�]E��!e#�/櫔�#F9�-מ�vƪ1V_�r�sp���"m��fdllA�nt|����ey0��J�.Q����Ph{
�z�'&?��jrs>�x<��>I�A�}]E��w@>��q4�|��@@��
$���g�͙�����ӌ=��4PTid�Q�@��	�����H`�X��!f�v!�kW�w�K��Y����a�D�j�c���?���̐�M�U��I�2бI)^|�h��A��+�p�}�<}�)��'�}�G$���N��z�|����+Y��9���0|�8��T,��N9{���reT^J�5�^��r�@���R�h[㶼)L��s�x�.89����
����c���f𪑏�>��]'��-b ��*S�y�>���F��b���(�cQ��. ��E��C��v������&��kb��.�9-�ё�~ϼt=5s��zF:w��]|��ؓV���dpJ3����)K����=�*?n_4'��l��.�Cw������cy���ڋA��W�d��� �/
�g���_}��������2�0��߀ 6�����HI��U��t���X���j�7�M1�[�,�ح�AT�;��FH�&ֽb��;�L@�}���^,�s��Q��y�0`f�l?�� dT�?�/h6�����s�| *,�:��a�26�3.���L�%�ug�y	7�K*��͏V��R�5��٬�;��U�!�mil��1�L�Eb�Z�ՍPw�-"6'e���TU���`<���G<
}&-���Nf�y;�/�$����W��+	����Ֆ����f~��?�������T�iy�s��
T:&|�=ȓ���>fi�a�O3Vu��q�i��k�C\N+�Dz������\��l�_��i�ӽ@����]�~�T����� ��h��8�����Ҩ�*b+��1iq�F&06�h��������;�%������xf́�� ��j<�$��$�N�L���x�� �8�kr]��4�1��D������M�ɇG��u7�#��|��[��h�?vM~�ڽMP�y\߮�'��c���ds�) ts|8u~�3f�E�����)�{L��]q��c�<�rr�P6*3&_���"�.p�)�C�$�F�,�|���t���z
��6\.��d��9r� N��HB�`U5�m#�������8����D��Rj>ۯ�!O�=��a���/�����mlٌ4?Z?�M���w�@woT������vHSK�Ɍ{,"a�A�vg���c�!�]�`�;�����&0��L�3.}�W����ndd
��h0X/���h�ED��Ͻ릛_U	���c�K�<_U�p|UBW��a�a}`:��K��W��7[�V����^$��|0��$!��	���<��)�:q��������(nR�n�����WȦ_��XXS]��2���6��E�? y�U����f"���.����i�N��2�j`�g"�n�XQ��m51��4�K�q�ӥP�M��|tN��t���\���i�!��Q;������!*V�JlO<��6��Y�,յm���uM>�����`�J߀��(��q�l烱�Fk�� �1S���y<�(F��E�v-O��p����x������^��A�ogmY=~���|��n���A��~ޑ/�
U�^W�����é��?60"&����Ӣ.�F�Cw|���T���?����;�0q~N5$A�ms>n�>�_^ҳ��>z~�n�,���� ��\�w��u�}�߀����`�(��O�����^?����n�;ؿ?�'�X$��Y	�e��JZ��^}T_p��=}���^2~���v�����$�o��ǽ�������~[9;�M�Q�Ԏ.%*�\��Yb/F�_��c)o��pضf����6�}���6.�0�}*��~Wfܝ�v�lo�t���ɾ`����(�񢷵S��p3�l���m�ϯr��h�� �y��fC���\!�r^���5Y��hwy� �q~�ʴ���*�����R~�J��n:��հ��oƔ�H�(�G���_��0�}���w�-?v��潥�U�b
Y�׫6��	.Ro���bj�&Ն	F�|l�? �	�Ŏ�@��G3��[�W��}J��la:�:Hج>wh�W��Y��t����o�`�̾�& ���`kz=\�:f�c`�=��4�M\�X"nxs4�^F��|J�ث?z-z选�[�	�}I�&���x��Fiw��[����lt�0�������t��k�7Mh��N0�Fvf�HJ��Y$��p��{w֗]��HJL�/"�ֵ�"�ˮ�e�Ky�@��5��}~���|��׋2o�� @NH e
���&}�?�0�\�b���S҄\:F�7v�yB���3'��v�������1�z:�f��؆~P��[4H���HPc3|�2�"9qY�c�����ib����Ag�x,6��j��?��x�@m4�qt����ԭ#
�!��^�C�fb)?
:a�]��@b	S�8� j��1a��pZ%2l`�z�{��
Z��8z��f�!���B��2rz��`;o�7f9m���C*����l��`Wmd�FE5lh���e4sSY+U��oc���b� �_[�@�h[�!�	b۴��25��##e�N������B�Fge���r)�T��Ơ���T/�F�ęr,}�V�!D��=�qJ�뤛�gh�����_K�3�Î�����cu�y}J����>���aw\�NL����H��l�d����WG��%20�3���q�	@�Ap��sUy����UU��#�Ke>~���������1���z}+ȏn�e�w����;���d�V�"i'_���Gf�����ˎ6[���g��k�0��<UUu@���O��k�B��
Lӻ%��\ȵ�)6�[�H�6��8�9*�P���k�.��%�
4�;��~���HǍ�����=鼷�Q�?�*)�"3��5�M$��j�1I���:Bl6��	�|�0fEj2+.R����qV&��(�)�mF_��p��O�,n����UD��b�~�Y���,3�a�a����Rj����9ao���j�	����5�:U�Xr�^_���
+�f����X�V�6�i��y@뉞���j������+���ĉp	[�^��M��@I�Pr�ˏ}��+&p���?6l��"��Ai���&���h�F����Itkd�ۘ�M�u�j��q���?��� ��^�{��s1`F[�SC��;��=(/bg��U���D�	�`�sqHIX�F�hUZ�hBy�/����l|n��9�zζ{��� ���� ���s�J����D��<Mg΃�K���*F�7�����=H��GZ�Qe�~�^�h���@A��Ѵ�=fz?�����5����Һ����O�����خ�6�^̈*]u��Ö+QG�@�(���g��sm�qB����ŢD0ᖋ��۶xՔa>�/Q���6�w��=~��i�t0G_^���ݞ�x�˴k%8�X���ña@���ǽ;��G��CG�	gr���
����xw�W���_�d&i���t����
������)
T�r'Eii�]H~�!�� ����F���E��e�3�Q��KTʚ�~kD4c>�z ~ ��f$V;�c������y���'(k�zo���EmD]���7ɿ̎n0|�@�!J�U���k4�@�c�9�Q\����Y�Ϩ{q.D6��y��N;�)?83ƽ��[���
k�[�� ٺ�n�l�Ā�ۦ�m��_8�-�Vg����4g?`�g��2��Rs}�×��d�TY4���&}��B�gm���}u9]X�
/��b�A5���m����l�o�%�)�MFj[�',���f�u'ry>�`v��������>1�Dj;'���Yǅ<�zp#�c	?��띾A} �nU��k����奥����ʱ�8�U����1���v�k�<ݻ��t,���Ɖ�����(�c��^���)�iS�r|�F�h���l?]��9&�ǝ��<�����@��fg;KPo��Wv�����ŅQc�])�W��d�4|}1;܃x����R�k���iI1w�Գ���0�}��|�Y7P��m�R����9h�A��MyCp�����x�7��5K����yq��Ud~k=;�=�+?�W��%������'mh�F+���=b�����)��_E"���l�s#JI8Z���z���z6�����=?��W=G^��5Xc"��� w=y�[��R��a�u;�7�<�P=�b)�p�w�]�l孫o����j;U��������~h.�{�^!sk���$���^#���K���Q��*��h꙼4}N�v%��� �*��-�]cc;s�Ę�W��N~�<L��&��p٥:�)���#;��2����4�~��E�h�#}� ���k~�>�%���S�bKK����R8��$go��\�����P���)��E�m` �W#r�*t�hٔ���7pSk��6ﵙ�^$#�'cG��k�5�;�ݝ��Aܙ�][.�G����0[7ꐼ+��*��xp�y��� w:���[����f�pS���i˜	� s&�Bg��|t�(%|eی�fh=YYM��AH�2�q���U:J��˽��oO��-vR��ˈ��zm����&��]�����.��L}�9��˞�ClH��纆']�x�a<�g���"����O^D���M(��,���U�x�fğa2����U�7�t���#���#r�@�`�����LHm�̓g�����D�֥���p�%W7+�
��`�N�uWX�q�QL+��o��΁^sNd��	g�y�iԲwr���^{4�s��<x�D�Eh�h����u��������G���Lx.%Bu�:�R~ԣ�s��ErfSO���+3q��yw�[nmZ�e��v�l�O��=��B�V�c�ϛ\�?����ڃ+H�9n�#��i�����C}�	H~ND7#���!J�Lm�ϵ���͍A��&���.� 䚩����,�S��M3�B�W����X�h�)�x�;Z���=l[�0�B,��
Qk�-���T�*m�v&X�����#a����]{�o��^���ˎM�.���R�^i��l~h��/o2�y�! F֊��a
�Rb��Y�uc�}Ǜ�"��z��n)��-�<��Y��ܪ�s-�K��2�����n xEh4~�+��f���+������1�|�9�!�M�׮Ȼ���Q]�`Ȱ������IS|� Hit#�����:>9��y�_U��;<m����z�w�y���W?��Ȑ���Ϸ���9��C��m�V&��\1��yOmBCk��IB��z�{Y��n�����<�N���ZY O����'W~q,�}H��j���3e~<2�x���e%T��u�E��	��9��!+��h���uӹ�̣;�_��#}�<ڲ�&��}T���ȭyE���ݱ�('��g�e _�kb�����h�j�s��L碍r��ϧ�(�1�y�|#�����*�y�vuy����f�Ҡ��(h@�����軣ʠ�?����� ��N��\U�_�&�o��Kc�a��0�j��Ң6��r��X�ɨl�j�?m��������{Me�nZ����:�܄��@�+?�� ��"��"�!G.�*Y���K�-z3��j��ܑ|΢3@y��w��p�Eq_n���m�D�׼2�Z{�4�����;��u+�Fkh>���R���:���V���V�f���8�˩W-�J�	��t�a�y		p�x�FAS'�\�4m���dT�=���+(�6�?5z�S�;L�WΛ�YR�z%D�7k��%� �{}��"6�0�@��t����m���'��x�=�-��5�p�����E�Nd�u�@*Ԍ�-o��Qk��^*���O�����F�6�R��8*J�Xܒ���bĝ3C(W�᷅�����}u��QhPW�+�@�mэ�*@��Jڄ�Ԗ�ԃ`��TM�o������)Q6���capIV?\��:` �7O�������2�几���Qq �����'"����'����`<O��Gʹ���M27.#5�j�\p��@��ք��&��WD��\/zu �ʥ�
�{Z3�ln��j(��c��O���R���n���e	�`-�M6q9����z��TXE�f��:�dq�+Q��ˑ���ʄW���Q~ǈ-��\�����6¥�!�{~�`��|�����t�� �k���(��>�Շ=	=<~b3wa4!`V���&0V'��i�Q��� �B�?�_Ʊ�ϟ}ښl9�N��:#�a�,E�dAdT�ז-��0��jQkݰ}�a58�.����;�fT��:C� [��g�Ѵ5v>��I��WJ�]�_gZ�q�����,�-j,�<�;� *ȯcp����6"�+tM�ًW�߻"�5��(������;�D���d���>F>�AY��=	��'cZ缒�/p������k|Ҟ��T���-�~�K��@�L�;@at���q��w{3s�Lpa�2��z��E�2t���h��fRtI�8n\��~4P�1�#˸+�0���n�J/JEW�6��/5�Vb�F�1u'�{���Ub���q�a�K�����X�?�r��\ƵH��G^�@{�>{����fO�0_�2�.��|�r��^jF�Ў��g�y�v�f�=�������ۋEN�*�ӵW!��V҄jc�u�B���q��������{��v,ٜ�r ��|.6=��U[48��u�*�.Z�\e�@��4V��������0Ꮢ�yRݹ�Ҷ�z�?�u�:qN�����l�@��D�_�����b@\�<>�D+�9Q��wM�����]�RT� �!AO���Hd����vK��h��Y�����������Jn��y�GV��[� ^�S��7Ltf��W��T_����V���Q�G�]N��KlL:����,�6�ט	g�僲�ށ�����9��b�����\�h��d��,,j�n����EQV-�瘽�m|p�s�:���Q^܃�Xݗ��k�;�i'J
��=�ix�,�佢;�9)4�U�>�E����ߛ�gs��~~�����P�ZZi%�����r�+yψ����Ph~�+z�&��- �k[����n�U���ToqYL�լ���T�΁�I��3������L�w��80�[��3K��	ٴ@��W���G\�h8j@�n��#Ɛ�WY��,��9�_�1��y�Ca���hQ94|ц޽i
e���@ktu����E��=�u�4(�Yx�Y���!ꁷ_�{��7��i���n�*
��51�^����y?j-xT�&Q�ܑ)?�"1�8���yM���nP�nW{��6��Ǵ�aڰ���ep;�UN�OW}�Lke��,y�+�:��/#R�8�a�c�뗍�KD	%#��$C��	vu�ͷob\*����b��Cv$�&MZ~t7VK��a�l�vL/6h�������D�k�3�:��łi���5����/����� >���sݱ
m������>�*R���9=��h.`G7l��� �rNۆŢ���-�5�G�SLJ��9����������$g�t�E��������`�c�r�r��ޔ�C1��c�.v~y�~*��Q "�Q�G���0Eֽ���X�^�J�bƽ��>�.��+壊#eDJ`�m!�3*�_�iLt3�Y�~����֖��CE��1������c!���ޥ�o�o�[�^�����6oA��o��a�^�wL��Ky�G�8�<�߭�h�'���R�iz`MP���11aޛi�Alh%+p�Iwh�"�{�1�%��]�~>@ɣVgP�̆@4���A g�F��}&�C���^�	������I\W�O�N V)���(�|N=Q"
�guV�'Ϟ�:�����n�w�2A��[!��_�mO2ƭ-3{�Є��((H������K4oXe?7 ���JgJ����j��G�^*%F�n�n[��-����0No��Cj�\��P�@������n��i>�"*�N)lk�ϼ�e�Zҍ(��q����8
̓Z�9���۹�ͭ8�  ���-S?��(��oJYXV3h1%1l��E�un$�f M��M�9�$:�����]��տ�>k]�����o������|��7����Ԕ��]?@�tcEG��]@��A��Ci{ *�ֵ��ۆ���V���aG�%=��YDvu�.s��jw��l�"i��^�H�®!�ed[R&�:s�~�@\I����-�Gg�̾�m����ś�r���]�փo�s�l?�Z��͞u;n�[��I���?�����l�hLE��m;
�Њ�pb���R=T����x����[���L��Hs3ۉ�	ơ�/K��w��Jv�w�c���s����kw�d_~T�;����r�1�#��yYO_FV�����R�c��;�nP�\7�)~ RʳQp������|��Bh?Ո{,	���ZY�T�Il�R�v�2`�6���$���w�t��*Z])���0>r� �`D` s��G� kǕ���t�����5G(�����K,�-���g5�,���`�����?��FFww�Ok�;(D����WO~�*�u�|_�[�^��~����J�֥Ŗ���EnQt�l�ؒ�Hn]��/�.wj��xոw\�B4Kohv���z�]�wU�	y}�pWꫡ�!�?ۋM�Mv&J�Fc�=h�*�۱r݈��!�]7t�3�E�X�y�&�n�z��[�)m�X���PBl:�wHA����6�9ˡfڲ3u\w��<�}�Gk����3����'Iu�G��Ū�>�Ҩt_�`�-�-����ܟ�1Z�2�D�t�Ūm��V+s��HTi,LO �3En���Lkh�7�I*a�Ы�4rߴ6�_�y���T�C��v�մ��?2�n����b���N���05Z��W���b�����̇A�,G�Hdb��<��s$(�UV�;��;N�QH��]�l���X���~���&4_��B�1��ڱE�c��Xu��I*���F�����8�m�(��S���讛f?(Ȍ���{ߖ���/v�Cy��>g.<�$�����C	�s=����k��ʍ���;�F��F��\�VR{���=&��ۃ3N��,�x�J��)�y�/�x<�C`}��_mw��^��'��{���
�Rh)>
���o�@M�|ĸ� ㍞G?����:��%��� /�i��Wi4Λ`_�v8v�S����;�yf�;5F߽#��8���C�X����AUb|�'�����M� �1k#ϻu2�Ď���_`?����2��}��¸=��s3�p>��3�X�X�x7���߀Tf�!p09��F�w��wۤ��3������v�{�.�N���T:����8�!s�&l�Z���
�(�>�Be�}7���I�����d�	$0b�7���{��zQY�hB$���~�b��\�:l�w����=č�_<زG���\�l5��:Gxx��`o�����To�����?P���\�=�o��|j,����-���8(K��B\뼯F�:�Y��������v_�6�4��	\?�N��Z��8�8���*��RO3�4�.����x�8����A��דu���Ie�kRQ�%]�ځ0Ғ�i{��#Q� {����`��<�+�4�ȑx#�v#�tnDH|��bv��6���ɮ�F4�"#��4��He���b��6��jI�/�Öj`���2�Yp�)Tt���6��qA�����}]����h~D=M�M�-/\�i+�L�����/!�s�������ﵽȩ���ӷ�:��ם��K˧�t�wg��/�p���9�F���$���G�� U��G*�)Q�����F�4�H�(�#����B|��/���ڤL�hs�]��с2�<�eYE����f�}61���r��b�Bz�ʁ$Ғ�Bo���7��A�1�OQ��R���'_��{?;�����'�S��xwT����=�U*�t|�y�>���;w�&Sчq
R�}�f3��s���R�E��\�W����[d*��~
(e=���m�Qݝ�ww:�hp��
�H�H�Te�R�����x�)Jg�ݣ�f��:�wF�z���������u�Fc� ��nT�~/>��䒪��S�2Y�n-
.@T�מ�S�ѯW�yIT�t4V��q���l��7���R
�DAܺr[R
���b$U!(YDʟ:P�2H 7V���8LBC7���^�[v�@��:�A��sc��ȣ��N)�;�TIO�T�;H(7�[�9>����f��V�q��j�����7����l�f�����U	����6:h�:�J$��N����6���)��G���1�GE�^谋��d(��R��]��똍=�lE����Uo����u�T��sP� )S��ԧ��I�*��w<�b|ǼME��w#z��U�a��<**�En\��OT,R�0�Qi��g.�A��I��8R'Í?�A�Vi](P�֩g�?b��;?���ԏ��
��m�|"R��6�cC������E�|Fk`1� �"��5�Z�֢c�x�j��F�ƛ4X����_��e���㑆�s���l#���?6	�N���"�sK)�r���5%*�.\�������q1X4�S��&{�=����M]@��|a����>�����K���^���;IQt��L�Ǐ�����4m�=��S�����T����|��&��kÑ�u�T�����o{x�6w-5/����ҡt�]9�n�B~&��b0�-,����g/&�}p~��l` �I�>9��9�JV��{�B&���|���z�?�.d
E@Cs�)`t3�Y`��d|*!6�:>蹡kN�zfR���Y��r7���f��\�%ڎ�sO��.k��@E�S�B@E��4�IƎk�Y_9�OWxG�R&)��KgA���v�j${:L/QJ�1��"c�?�F$�ɺ �T��M8E�3L��i�[U�Z��0�F��2sT"r|_�tg=w�����ď{=ە4kK	���7�U�zA큪Ǝ{|_�r:�/�'� ����'��]�W��IC~�3],�@[���{<-С¤#����S�	��u"o��Lw�1�>����?��d�R
*Q���Pe<��QH��l�XF�h�����03jtbN�3JH���E�&�N�����ρp�w'}��ZNB�kU)`K�;z.���A���v�O|�O�q�=�K]*���>�e�eMi��G8C����nk�Y�q�&&X���4�y����� ���0>,^R�رǝ��#Ď`���)Ad�;ϊ$rJ\�R� �6�._�ZS���37H��#1�$��
�,ҿ�T	�dB�Xm/P���s'\���M���텾��?��3�xR
yI���>Vu�p�9u_>lW����Bȸ�A�t-m�0I����>��S�E����ظ�^�6�l�S�Yh���t�c3�vy�YNvvSA�C��E��i��Zhi�rB�j߳�}@�G�B��G5IE�ܣ\�#�i?T��%���^CD̹>I�������o�9�}����u>�̍�����/,3"B\�:%/4������-A
�CcZ+%��?L��ǳ�K��Q{��v �}�Q]����F<-���7�'�b!1wA�-�F+�	�$=���I�U!�/6�)�y���Yo0~�һ�xG�u���W���y���yݕ�Mi?H���R�U�C"��İȎk ��P4���-�S]�z��ޘ��i����8F8�VQ��r��tuq �x<��{CڨY�A*�*�}'�5Y�� 坸��ڣ0�^OU�漼�w��v�_<���w��q������^Ǽ4a7	���c�ip�������1�=G�$1.�v
y�D*J6�c�I=j
X�<M�T,mS_h�]�͢��?�!���D���nH%�M3�g�V�% �=��:I��{z=�ힱ�g�k�4/m�ὶ��5Ǎx|���yc�m���d�!� ��b6�>��8#MD��7�.�.������U�c����KUE�)^�[�3�riTG	�(�^O�!����-��^�Bm��F�G��F�aix��߷��ukwRHч��8�E�7k`�s�#~���p\קCޞ��#�����ee��W�D��<��V�y6���U�~=��5R��	��Љ�2�:�����?tg����k����z~�@�zU��ՙ�ACG�����.��dtgX��i�v��rikmZm.:��Gm����W��?�/Y�u�|��>N��J9����KT�(�h_t����}c
��61�MB�}"��	TN���ߔ��_�����[K�m�zA�2nC�LnޝL��pA���U/���}�s\W)L��W��!���ނ/�S�T9rHݺ;s|U�GW��@S���}}��N�d�(öa%�T��?.�2�\��6N/"�sX��l�੒���)�������c�i�Ru���wܠ;ޟ	�����ö2��^A���J�ꕩ����M c��FMs� &���Kez��񺛂V֝W[L��3��on����A�iAA�Z�ڍ���(���chf�$KƗ !�	`����D�wY=@dF��'�Rk#��mi�+u����C�=�%�����Xڽ������l������>���7�l��� '�����m��%���ZUɢZ�ǡ��6��(�i�X��� ���;Zd	Xu�@'PP5��|�r���X��%t��ye�&>8�Zc�K�b��*K
/A�+V{ؘ/��v�.�n??D=����������,���=thʲY诿�g�wӇ�M� _m�	k���]�c�2*z���:0��P���v�]=�=��e��~�<������؃�zG��.Hi8�w�	ZPv�&g#�WV{㞎��lT�?x���6"���K�_��7R6����_j�ũD�t�̏�="hK�ۄ����j�^^��(L�����D{%̶�	Y��-�@�l�;>�^9/U�6_]��T��]���EfDq�A�*�e�Q�����]��l�$
!d� �����pT$n� ��t-s�AC}�\8���}= �π٘��� �>F���C���4�j�@����q_г0��Xx�����fUA�2k;��U�j�.�-)U�"jb+ �[ec��'1����? #��ٙۧ6���=;�d��K��%4��]�h8���s���i��3�6����k�ю*�.ږ	,j��y�����46g6l���>������^{�?�[��0��+'�hY
|��Ϲ?Z�>I�g �G7vOZN�議N���v}$��=��[A��U���zyߩ��Ƥ�r�͚���(�*vt�"�1�N
%ڏYk�\�SV�"��Wvk�������|+��c�;���6���~5U>��L�*��4aclP��Z�|��7�P�J:dA��ƣ�u	Z�t}i�߸�H�;
Ft�{@�� ޵�B�&JBL΃L@e>�{ߩ��o(>!�/�����$����h	�iFW� ����{����e�����݁��H�!y�ڭ(P^����ǽK@&��Tj%R�4��v�w=�;��Qd!����h'=��2�{_����>�z�,L�/��������aJ�"�;�v�B��q�����ij�<fE{�A�9�M�]�iC��D��q
इ�����	w?Y Ȥ <Z��j}W [K���⡩��@���Oer�R;a��dg^�}�_d�PJ���/ކ�j⁯�*��] �E��v��N>9����Ǜ�	���������*�'$�A��M}�((X(k�:Z���O�Ime��
 l� 0D/	poҐ'���S��(�\9����T���5TQ8����w��)|z}����4�?z;��A��a���vt�*.2����Ƃ�Fe����V 3�8�~���N����]�L� ЈksXd�$�������y��in-�ȴzA�`�s(�̣�rw%C�������2�H-cj�cr��-�W��i��_8�����O���g�6T��M��!M�:��Qf�#: =j�@.�>9��@� ����[aK5l��� 6��������:&d����5i���+B�[i�=�*n!�{����:���Gʸ�e!����;8�e�������rר_�������K��;Zo�QEtN���O�H��A�f"l2ɯ3(B$���	�qDfZ�v;>`)5[C,�"v��4t��;%��h����v�d���*��R�	�NA�^�^�j�,>#4s��Ћ�1wjib�Gpˣ�����F)76g����\�n�F���fV�}u��GM�P�)�)R����[�MJ�HCD�ų��fM���zB����vc�|؉tE��D({4�mMd�3 �e�UN�}�j(�~=<���T�~�Ka����p�9���Y���g�6��z�/��VoV|��'�7�Se��Wb
�`��4	�h]ʏ1�,XD�`�4�ċ!���^�Y����y���IN%�q�z-���")��w���Lb"��%m?�h$<H��}2�ߞ�֥3��qW�iG@�_��:j�p.��1fX�nb,(
��l�58�l�@�Ҟ�j�se������gMj��zm7,�v�A��*�w;�(�Nc��O�Ղ��F������Q����O'z@�]E�� (��q:>p}�ۏH]���H�|�A���3��z��^��U�X�]i�"�QGN"#�0�|��H��	ۙ�^�su�E6A�u���9]���߻�e}p_�ӑ���z@f���[b�Z�0O��}Nm�5��j�9����$����aT�j��Ɯ���M\t����='�>&Uh~���Z��D���H�;Ʃ+����ո|���ݪ����QQ1��}+�}3�H��f
A�5DZ$~&�X�$� ��vfUY�I[��\�!��#w F{|lx��X'=.M��#����l|��u���g�	���-��C��+]����X}k��O�(�j�5��i�|�f?�<�XtZ����E��1씅C#kQ~<ʚTTZ4�jJ(��v{���	t�z����ޫ�xJ�0w���6o#j�O�Ϊ���es��-���C�(��P��Jw;�n�f�iX�~�i��H>����x_����z��g!��q�D�dx[�^n��QSʗ�	�xq�/ MG�t�EM��D>��A��W��I�sQ��c���Ó���C���sO�QjdF 2��)j>�;dfÑ�1C\0p�ne�Uo.T/����/]��ή���Y�+E`�7��X؊�Y�5��[X�2��W��Q@��Dr<���W�k�1)���@��t6G�ƿ%Ho��Hjx��R�
m�h��W�q��Gm�2g�l�w�򇢽�,b#�l�GFp�O���y��i
���Z�]�RR���lb�S�*)�Ɍ�o��˸��bͪ!׭w��`B�C�W��f�x���x6����X�9F��;��C��¤~�ʴ&�^[��^2�g�D6f�����>��i"����n���/�X��U���?U�su���=V�lh�R�Io��v�&��V���UCG�>�(a�����gc`M1�d��0҂���آ�%� `�6@�[�a�� Ҕ�Z�!�߻�� ��|m4X�� !��+�9B��Y�<��r �3ߺWwJ��Ǻ�{ɩ_��ύ��\�k��F�sw�g `��Q�r�J�oZ+Ҥ�E��ω� ���X\�{�hL��َtoN�&�� &�tQ��C�U�g�:hKs��{���xy���˫��!B�	.��I���_X�GK�x>Bšu�ɣ�96��YӴ������(�]Τh���(�s(��{��8�)KG5���>[ً�b���?��M�T9��|. k�!�Ge�Ch��Kց8t��4�(��2Tɉ�|ܗ4�U�-���#���>;Ez2��eq��_R�ԍ�2Xb��xGS�Ƴ��_H�/1�ʩ�0�I9�&QdT�S��؟��u%Rk ����)&�(2��)s�Z��죡?Q��L��G���n���A��A$U2<�Q5� N��:���,4�Z<D7�.Q��NZ2�a��0Eȑ�O~jj�7�����2P�1�ܚl���h;y�P7�gF���NZ�����D!���xs6'�|jC��r�L��Do?��ڽ1�S���BB������R��A1?'��c*m=",�q��&�
Y�ƈ��CۇE^�����=M&�`q6(����~o��+
j���M�^� e�'�3�/'zhm"�Ӿ�>�`~/�F����T2T6���M�У�|�1��w�2ϗ����u�sSE'�xC+SG���h� �����j��_rȃ�m,���Q�5��b�Q��V�$��(�A�vd���a�nR�;ĭr�S]����&�H��g��=4�{�����>�����Mu��y��?g��p�/��,��t�*L��;_ut���r���p�s�p߇��V|�
	�f�����U�(��؟�(��TYN;`�TwU�z,;��j���/��@�C��>�%� �r��_�AJ�������(�E O��]��=�m���t�j�w
����z/t�DQ��eS���O �v���ž3���F��m J)f����i)�[��ud�Ba3�.Awm]8�+Z�;�N���@ߓ���*%|���x
��i�PK?c|ڀo�� �6,�-�?����o�(,��k+Z<��eFs����k����W"~�R�zm�w9�����{��o�"��a�Q��K��(��S$�(�;CRw����fgi/@�|�^P�Q��>���#�`z;�����LwǝZ��|>��#"q&PC�J5㻸���G��ܒ�ozN�)l�i56M��Tuɭ[�v7��|�;Nt���r���[{Λuވ�~׏��#�P�cKͦ;�nW[a�gbi�=����!K�"�oCx�?0O����7P��-�d�����ԣ�hJшU@�Ds.�[�����^�*�P{�Q:ؿ�  ��2��u:���J���tg����]�	#b#,�)�����K���V;�摎��Mv�5N%�ݦ��m 7�B�cf�=-��@q*۲h��ڢb��0nw������A�I�(@��S�������%�w5n��b�.���,��4:���`����8a/!w�Z0�!��:�i�?�0�F������/�q��<	(�)$!P��U�"{Z8�4��/.~��@��9:]ؾ����蔀cX�L&�)kqO1����o:)�&�{U���Rz5��E��7zʏ6�B�v#�R���ZO�LX:�څ�t�MjB�aj��Jl�@���#T�#��C=�Y��Q��g��g_B�{�[�F:Eɍ�������@7�lm@kB����&�¶3�=�*�f��j?B�>�CAOyc!����\���hL)r�R�n(c��"���F�Ʈ��2��%�|��8�*�Ӱ�^9�2:�̻�J9n1��:���B�iU�n#�&`�0M
z� FD����r���_.�ƙPB{V�"�����}�Gb9E��~�ޖ�v�I�yhc�Ɲ��~#��[Dr-�ac5]-�����@9�⫐���|�g��m�!c�	�q~-�ެ͸�`Ӿ+��i(	���!}5|h��T�n����ث�U�
j$B>Е]��KCL�B�	J��KU֥X���1B���Ԅ7�ߚ��3��.��O������0A8�U����EC?)�w����j8`57��0�=����6�
�����%A�#��M]n����f'��h!�uY��6�j��҅O����l��j�]�K�^��m���+%H�Z �3�ϫ�L�)���tnÒ��6{��<��M�g�[^����Þa4�*i?u}�n.��ޖ͊�
MH�|�$�O�+-���G�\W�h�	���>�eNz4�NW�i����'.�r<�З����F��\͈�����ZtW�F�����!���ՇV�0���]�~�_l�[��4���W^Y)�&���+�p�+G'�wͨ' �5F���*�X�pQ�����ᴏ]`���G��x]=a�G0.:�~l���v���H7CoW�z@ ��M�~�v o�?���TZ�����������J�T��r>B>�����Bj����I.�ƽ�z���	�C+֖)�(8��m�����:i)��wE�:O@����^	Q��%݃���i4����uvgb�G��|io}��*���t���py���~�MƫM�&G�����}��߈R�nX��ZH�Q��o��g�z��]����*5m��>��|𱚓QA
�r7�:�
�PeΘ��;c��yJ�w���;�,�i�T�Ih<��8��T�����h�[�xEv���*��C��<:c y�n(��kw����ʷb�xBv!(!Ǡ���s��e0!*>��Ѣ?����>��zu)�Iq��A���JC�?����f�G�U2Fk����*�@BG�f-
8�ՙ$�
�@�࿙��~�Dr+�rs�&����@���C��=�'��K��dQѬ�Ԝ�d\G2�ܾ��
��hnn�gY��/Z.c2��\DD���z�����ә�woRP��8T&cѭAg[�>�ָ���3\�O�[�,����'�ܩ7��'�]W�.����4�=��=c��L������U�S��]	���o��:4a����ps�ҝ����r��� ���-WQ��W�"�a�0P�	�[��ݷ@��3�N:Q���}�2(Е"`�ZA�"�"F��i�?�K���~��k(�c�g[+�5ik��{Pr�C_!Xy7�x���M�>�:�J8��xg�Ť��I��'-]��n�q�}kD=�B*�(�p�(霆�kn�`3oL�a�/_��3�X�=և�1n,M�a��ttI��!�I�t��?�K��G(d���T����`�9J�,�A6٩�u\�׌�kl��ݗ���m�>˸^�A�1A8 `;�U���#BoH�FGO5~±���,�QOd��|#�(��)Zp�̍�}�� H�f��#i�P�վω6����bvָ+�s^���)��e��/?���a\΅I#�{�!�%!R��*O�&�K��qL�� ��+�� �����PE� �#HjM:�
B�۱��<��u�V�wJ�-E|�		��z�d�x��Ϸ�X)"^x�G����d;���G[(�'*�aDM��Po�zf�r��QX���c/��ՙ���cI�k
�إQ�R4� �!;�<�����	]�8w���v�θ'��׉���Z��T�u#U��-�Z���J���r���6x�H�L4�DU���

JN&����Ɋ��/V�W�Yh�n:�x��m���)i�E�C��G��GT��}#U�%s����Y{�(Xm�{�F!��F
i�3�&��LS/�Nc
Ky ��q�����J�� �ګn�W�tn�N�nԻ�~X���0�lRAtG(LuE�;��cМ1vf4Q`�����F�2�/20�Oy�s��Z�Of���m�?�b�a�רy��Wݷ��6�p=U?��̹���y��l%˾x
�\�l�z�!��|\��[�G_��y�3X_��KYoZіg�+\�-��}�L��W��7�=��z�'���o���L�Q�`�xw����B��=��Cc�B�63���C�1sA�|��v?�1����_z۟�񙣧��=[}�us�"��-q
C��ݫ�CǗX8�*������R��.��]���0�`#"4U�t)5���4Ǘ+ߐ�Y��LNr�) �N=㺶.sC	z���'�ߧ>k(`���.)K6������|�K���ц��6�9��H��;
�}�q��}b�]a�J?��I���c����9Q�T��3�-�tN��3�:9�e��.^��7������� u>!�z������wF~(�9@�rOrR�例����oq�ٵ�v;��5���z����*}FثZ]���bQ��6�\�A^Rb��=&B9���]�x�:� 5��r�#��c�B���D���ܾљ>��_����*��*�p� �j�~�R�}#o�EuVG�.��{�Y��7�p\�
���h��#��j5�9��Y����1n��â^~^w����'����jۼ����z��D���q���k'S�G�sW8aL�d	d�0��E�^��/!a����5��V�M��V�<�3�;iz�_����(M�]= SK�U���bmQ�F��Md�Z���@*^�Ԍ�FaW=0�1��o���§k�{]��ñ3~I1��j�.w?�����~C�Eِ@��ek~a�9��mv
gM2S���:�����/��qEY	�s\*ƶ�dv��sǼ�^���a]Q�,�'G(��$B�X�]B{g��E�>d9�n '��Ð�2��k2�MB���@O��<{�c�3�<���<�AmY�ku�2h�3Q�b���/��{>A	K 䏆�z���������Q��9�eܟNmY���hZQݥ��6-��n_����!&��*����ӄ o�����G����Hb/����>����>�,�2�h������s�Q\eW���f����~X�l�ei=��IHXpK�M�1zC�D�H�6�89��ǍrV�S����9Q�;��l]�q8"6�7G͝(9~,����e���=�{���f��M&�U��A���g�9'�b>��
Ao&�c;O/M ��ú	��T�qLn��4��~uNݦ�(��G�S5P��,�=&�Y`�&'Q{�ԑЏ#Ao�t`���T��3�p�;������fz�֤�a�gщ�Lp-��9%�om#7��갽]��ѡ뷾�[�Blj��߬؁y�Ka��G��iC��Ɓ����2������r�we� xo銪�D�������j�ԗf�g5{����?�@b:j�<���#ȸ`[٢x@-��1��Ǣ�f�����w5��	K#��J���L>Mft���y��՗����Zi�[�MGͲ�tO8���݁�4���V"ĥ]E�U6��x��ir�5��:(�����W5(��Yy#�u����B}�ժ�[4��G�B���C�`�|.�bL��Fl��w_�m��o�A�q(x5O�u3]w��V+���b3��(OPM�vQ@'O��߯�v7W���#�}�����>oS��)$>�I�.�r/�PC�$�\� e�`��`e��x�CX�X���s���E�J<�t�����ڕ��9Ju
��9���Z�T����u}��IYn�fg"V�����D2Z��'�#��:*=�Qe�Z鰱Z�RcVT՗S���K=����ϻ�x$���CT�&t����"o�k��q���ՉK{`�Ø�W��)���hN)a��H������@�&bm:�£�?p&`����0�B?�:)�
�>�K�$mM<~���Z���S�-@�G�K3\%���q���u81�A"ML��:�tj�t�QYrҾ�Ͽ�9�L�V���2׫������cי2ގzՉ��W�E/�e��f�P�\]�������2a�ؽ��d�8�=���W���os8^h�_sHG1n���p���(�D:�)�s���UԆt:�!��J�k�j���1*o����!3�?)@r'���O�߰q�������>K�g�<X�㌻�����ſ?��Ñ��8�5����J2���7��"Ŀ�K��`�or�p���0�Cl�+���q勄�9�v�����2���ܶ��.���O<TjSZ�)`Xw�C��2:R�5�&=vn�J���X�Y܋��>>��f@	4\愿;�t��B��ۉ��C9��į��X}$	�|�6���ۡF��vp$��>x�����v��`��J�pL\"��@��^X^>��Ɨ�M�o���G�n<L�&��l��;��E��ߙd,��ƦB����y6�ЃF�j��qͰZ��!�c��E��D.��i�Ym����9���?H��oî�(O����h%�s=�`�9���S�9�Q& �Q�����@y��>�c��5���J/�=����?��l�A��'�3�#�O���������?'��V\�kA�W���e������`�)x�����f-����ZVD�XdJ�ϖ\��ٖP���E�K�|��p���6�0����F�):9()m�A!����Ga�-�}aF;�Y����q͋tu��1\ۈ4 ���=H0gȤ����Y�3��ݨs��]p���=�>un�l��:�B}y6;��o�\qH�~�m�x� ⻦��n�
&<It����ߎc�UIщּ_�����(�D�y���D�4�:s�]T ��x9�at|w�(E��n-�(LF�=�����4NA3��(����Mu�-t��K���#]{��NmZs�K��]{]�Ⱥ�zy��(#��	'jGd\����|���됳����mL����|Pl���TD^���]P�:�5�����my�[������d�A���;����Tz��'�����囦���|���Q�gA�~��+�%y�Ҳl�k���yJ�RH���M%��1��kb�nFH�����K�E���K����dfv�#��%!��G��J�@�A���tnU9�B�A�G�p���x'	4w�`g��yI5k \�[��K���|�9� �ܾ�_����w�y�?E�-B�h����(HU/@w��V"���a18������{sq�/ۀT����>ǩes}�f���G4+#+�b�~��Æc��8����G�RWe�/J�?���^gҳEs����1 {�K�0�o`-�����7Π��W�@�1̞�p���+��2ТK�VB&�M��:��h��Ss�0%{�o[��u?�����"ѝ�>qT�h?d�|6�s88S���Aa<��؍I�z�j��3�.�"�T���#��� t�*r�u}T%�,rר�sGG!hWP����K����EI5u��;�B��W�((��^k �]�.ɤM����)��]
6D���V����h�i�JT@�ց��5���TD	G(�VJ�K���3���Z�$d�o��ԒQ�e������	�*�alP^�;Le!ga��8q���i��
sM\����`Zp�������4�ug�[{1�]�/�N�ۊ�P�уk�d�������Ӯ͆7���ㆧ�����(�s���܁� ������G�qg�T�[����"N��,a��Tq�֣Z�稣�5T.��>�b�W��� �B���(���I��@?4 Y��̪L������he+/}4 8�{�2�04iN[�JR�a�-�"צ�p>z~��@S�_&���w���M�ߨ���g��x�8�j�4��&�&wǇ�kE��H�_��_���T�fAv)�D_��h��$����,L/�pS���������>���{��	�xQ:3ʼ��G;r�6�}l��.�f��y�;YS����A���R�|�J�fu�FTUɫ�u�o�_�o:��2Ne;�NOT(�=2��Bո*�<����~�Ry�8�kFTT�;E�Q@Zw�y��:c��Ζ~��D#y�I��J�{pq�OT�[��ra�o�~_��wR�P)G�0"	�A����xZ�m��N�_�Z7"|�c���-�&�(!5nQ�j�^��ﾁ�ƟQ������������P���w�<�}��%1�-�ur����լ�����Z��{WdW�!lG/��;>��pXΈe��8�F��4�:��+�C�}n�qn�D]4xYo!��	;�Z�<�uj<�6�Ӊ�K��p2��J���Cn�=������j��Ր�|��y���/����r��F��2�n������~���D�h��)7�;�d9{��@� _*R���j�^ ���EV��y�Ʌ@� E����1�rtb#s��m)�~�4R��ߟ$A�)��O����=�]�M���D��0-��r�����	с#E-�P\AY-5t��6�6��y��wq>����R�<��2����j�A�W�&�sm�I�\��￥�@�ܟl�T������@�ﰤ~q�#;�3r
���a���ǊZ�&�(�X�vE!��7%�A���؛DË�D�DY����!
�pW�h���;|���KB{�c��P�����v��o�aW��]ӏ�݇	fV�^]�@,��=*����ZK>0��r��s��vk_�^7&�;�W9��?X�"[s.BV�,h2���Qe��<�5#� �����K��5 �EՈ��hN`9Iֻ���`d�zM��XV~�u�����X���B/-##�J���n�ϗ`�_=��s)h��&�Ix�~�a&M�SE;,���v��Fi���2;Y2`v��Ū0�7.�Z��溡�ئߍ��C�YI�s�]��O�T�]�_2`���Y�K�~�K�)�㠇Ej��{�5�Yq~��]J�݁|3F�.�Η]��%I�W��z��/��:�P��CmA� B��GG�g�ݘrh�w���C�^�-X�y�ٹ���]~��<���:`�72p�(�h��@،G5ۇY��y���BS*B��h�G��%Y�%�s��@䪐E�~�=�c�U6"���f��<&�����?o���u	�b�ɉ����A.�^��@}��l0�����Z�=�A��쇝��/��o�@� ��hMz[��ma�7\쥜#e4����wp�B�8�qvng`3�#h�]O��ն˫���@}�(�Y�~���Ll��[#�����}k�����<�7JTd� F�cޯ?T���B��ެM�9��� �E��p�׃jW�k�k�]�/�Gى�=T�20$.C��Yu+|�%�$xk��&��~���zI��p�w}��I!p$E)���*C�
���b�
�owcg�{��|AU��h��?�l.[T�l��]ǵ��P[����+��a���:l&��F��1H���s��
�h	��i��\���R��=�@�*K@x:28�B�I�<?��=V��>�Sc��� 4�gZe��
��N��d�=u��v�F�M���@Ē�?�:���x�8"d��@I����Ta%��tv��Z5$W?�&%J*���󨖣	��2��R�%NTy��PFߠud���c`F��� kK��(���"�%�x����`��u���9�?j�ͯ{흗�>N)W�	����}���u���،e!�Ѷ�g����l�����-������V$n��E���M%�Ov�m�@u�2�2Q>0���'F�����8i�z�ñq�IYNŹoC���KZ�����Px:���&��c+`!Z����^P̋huׅi6k���['�u����x`KW���s��T�c��8\6,�.Ҧ��;:~
�Z�|ն�ϋ=C��}ܯ��n�ʰ)ē@��q����|����I��2�Vq�P�cY�#�;�muW^��`����~]�s�CA9[�*�.�]�b�Д�Y�i��w����]��x4��m>��Oń�� +�.H&L6TX���o�Qi��ܟ�F�T2_�dw�$���L�=�}h����Wǻ��/��֮��a����|n�%v��7�9X�q�#-��kygY<�ڄJP͸@�]�6N����k*���w�,�� '�ٵ�.m4���d�pP���3�Y�xS�>���G<�3��Η�ϧ��q��LŌ1g�V^xKx�sXE�r���ȥ�l܏/��J��2LJ����;�^~ �����7LKθ"nH���h��w��/���MI�L�GRr��@1�l���Ѩ.�'�ڇ}t��q�!SUp�^G%�n��Xm�3.BM��5�8�����0ެT�cj��0�Y��A�b���xn�}�`&VHB�9�����%�.�c�z#�eO��Z�~o ���=�ojB&�q�DbZQ�h��~C���G�f�6|�P�� �^�8dY��x�ݖFg�>�-�	�Qӣ5�V�{�w��$ou|��{��8��;���I|���h�(�n�-f��!�ZY�6ma0+���^Q%M�!v��lw�- ��*'�[��h֡oBY��Z�Y̈́������	̑�}%+��xZr�~���� >X���T�Q��t��zxw��&4W��[����o��U���yn�@Kk�N"�ƭ�|
G%2�s]U;�C}6��D%�̨�����/���(bϞ9=Jw$x�<�-��Sغ?���;Uy��<$=tI������ƹ�6��S��sX�o�&Un<<y�ܲ�&�/�O���7��q�����J���p��`���Cc��ߢ&�uI���qbv������"��x���ï�q��5��2�����"D���٫��!wT�V.���S�U�E��wdt�f�}��Y�m�ma"<hY����ɷ �}y�]��R�i�����p��4�z�^Z�� �"�Y��ȏQ��JC�$"i,
3^-��(�ٕ���w�*
oT����f'�.Z0�",��P��`afj���k���9ȻceEkj"��"=����ᐈnrJ:eKC�(�uc��W6C�y��!u`Pͫ�W����4�R$�<E�h���t\5����N�8��OE�xG}E������Ӄ�[��Ѩ��m቙��'��8~�@i�0��JZ(����]_[��RЦ��{��y�6��51�d��$���T�צ�V��6���I �=�f��7+B�Ph�nУ�b�=���1���{��X�K$����������'�CL5fT/��:��v\|�#����]�����5���Ֆx���rcBV�B��m���xE�@�����Zϳ�ȴ~;~�hr������[�Ԏ񃾏9i�+|,��q�d^Bi]W��b�S��6R�$땃�t-J�hMU�_4g���?�*w#9@dv�E�!S���v�i������秂�B���ί`��|'?ů�ӫ������Q�P�
��b�7TAk����)���qA!�&;���P}1�T�]Mƭ��Qb/&�>Q�{2����i�1h��ڝ���/��K��v'�#'��u�����("��+��,��;�x��{�;�w^��B4���[���J8"�&R|��p�'N��zޡ�Ey��Ɉ����
��
Њ����K��i�s,/wǄ�r_�c������;�5��Jù�n��T�(�k�c�n�s������0aO`
}/AG�NŘ��g>@m�n �H�˻h��"b��b�9^��{��]���_ڣ�I�U���]��5T�/uUvl��(�@��@�<�	��&~2�5S��hQ-N�]�l)����\�����
�(J�"U��.$4�����v܇)>�g?o]�gB����@�/B�>q�� :���렍:�1�'C�6ny��?�B='���w�8�� L��(iINI�;��Gٹ��w����΂���T+B:�0���ԑ�&'�.o2���h�0����C0��9�k�x�v�/���F��x-��Tmu�[g^�<�Q�'Va
u��!�aC�Nye��T(�2�u_��TW��d��d0����������E�CF������$��#�'��ѐN�_���J`������ѕJ�v�}����hU���Z}i�C���dT�����llN*�4�gf���W�R�����@EO<
��P�?�>����<�JW���8����Cg�Z)�vЦkr������rD2�f�N�/S��]a>�Ϡ����Ӧ�n�X���-���m�j7�����^��Ҍ�Gb�"B%�(Ős;X\2߈�OUA��,�9sT��=XTu�v<��ky�Y���Ƚ-����ܡuWTG8dn��IY��7�.njd	�޻�G�퟾I�:��u@U�+�Mb���<4��s��y�=���y� �)%M6arèZ�E� �	�~�I�?�@��7��~��~��q���W]�wM<Hb7��r�]�x�\ю��,��vC1�<��� <C�F�7鸽��a����#�IM�t �#ܛ��*�S��v1���;���/}<M���~�����ٓv,�����VM��7���݊�g_/�c]�=�ڡFE�R!��
���#u��J8fcޤ��~(R.��J�I�X
�z�)H.	!=���11���K�EcA�FidU��i�s��_��w���d|y� c��"T�+�� �Fp/�F'�
ʍ(�8��	�n46�Y7�a�r?�h�P����9C���ꕜR�D���A�zݸ^:C�-�-����f����,�:�D7�mH�*rN`|}��8��}G銹�� ����7W�{�U�)�`� �?�K������#�tI�K28�vb~-W+?$UG��:�F��u��S�B�;�W�SR�@NiKh�s�6��I�� +:�& �*j&�ĈM\��D@��뷎��|�ꬠX�A^3�=�=��ao��X�V������!F	��{����o�~^����箻H�HM8���R�o��qN`�ju��.=��ؙx64E���By9̈��Z�eQ%����ٮ`h�(�[ᘷ$
ݿ�D�2��>kC��+�9\��W+�����;� �����\ 衱9_s�7u�B0�a78)��		�\���9@�O��dД��w�s�qğʍ��LI#A/�^���Jf3�j �� �tA�Q²�x���j��ٲ_&��j߆��T?lz��Ǣ�����WK��u����,��٤5�v�*�f��r�2����~׃V
��.��y[d���N�)�rׄ��:��ޖX!G�e��!^��gc�� ��������0��ۧ8bt �Namv��~w�R�$���P&��9pި^��T�L#�hY��ͣ�e����%@��р�y�;���lz���w��;q9XE�g��c[;&��(�5U������;�y~8_��bJ��ã��,�]A ��=��SJ��
mV~�a���>Z��� ��&P�K�b7����:/�Hs�~F���_�я������@��Y��Ƴ��mD&����Vq�k.@�H`�ZA�Jw�;���|߽~�7�w#��;ɥ�G.q�(�0Ym�Cr�w/8�k�-�h�)~&�h6c0�c*\57�us�`�.�amD}�1��a�s��R����%7MHj�}��$��e���ф�׽Dcۥ=�Mv��O��:��DYy��bS�8���J� �����좻ߗ���{G�31���-����SP�S@�;6+��/6k�l�]f���܁)�"�O|ys���<+S�y��D	���F-�����_�Cƌ�z��i����+��F�}���ۙ/����y�)&�(�D h��r4t *>_���!z�_?"����k���~���U��r�k�fs��j�]�E��q��hD$�]+X?�
���/7�]��je��/�l��M9�<9Ti���`����S���ܡ��k�Dc��
�[�R8�Y��A��BٻO�Rs$�g�:���R�f 8�c�!��>~���7��3�8F�v����^�T�6٬֐*M�R���l�f�* �%Q�
�}�$�?����)�Ae���A��)�rR��6���Z���(� �9��&,˶q�C�٨��.�NVc�W�lۊb�37�J=F|�u��Օ���T2�C�mj���n,�(�N�o����t��c;�|���Z���(�ދH���V��t��>ҳ����{ *EuO�#����]F�v{wN��g|�S��Ϊ.���5t�^���m_+��������:'���,�s����������������֩�ڍގ�YZ�ѷܩ���� �u���5v�#�8�uAn޳TK��8��L"�ƞa��1\��Ib0���*V�sޢ����>t�#=q����fFa�v��Q_Й&*���x��w;p��ߊ簓ͺN5d���G�Ʒ5��I��<{n�Z�6pQ��)�Tqetf�U�g���p.xiC��X��DoxVq�iz�m`���,��z���q�e�sIBjV��E��wTOs��j�r �5e�z�q\B���A����˘���_l�%SjZ�	��$�R����[�jNj���"Eqxߋ��>��E�[(2T£�E�� jؕ�����g�������H��������9�s��ߟ{�]��??�<~4�F�{�ǣ3e\C�UqN?ҿ��v�ѢOh�Ih���	�faT9w�J�7��@r�9ݨ��Ì�<k�����R�2�.`�==�(�uE̎J\"e�2�\�s����rS��Wޏe�zA�����G���<ENC�x�l�ή����N����y1i��G4��N/��Ψ>�$�j%��Q�Q�2R&�'��F��L�����!6������Ѕ���������̜3'֫l��ڽ8i����Ȥ "�ˉ�ΤqKe�{YAo�r����t����Н���cw7FO����و�RM��H�l�s/�NC��,L"����^���STQ��� �0@�t'�Qh����o�2Nj)�<R'��&�0=��o��e�D�d�8oY�a�~_[�2��s��7�,�w�S��7%}��}ɋ�fRDs*�D�l�k����\��*1jC#W��V��r"`u��{���)C�>n�@W�q�����Nc��|��u����z_\�{�S��l��}�_�3���
�i�L�{>6;�z�lB�E�(#E�s�t�ff��P��*���ؾ)���F�Z�>ٗ��Խ��/g�1!�άr �f�{Ǘ�4e��E� �A�d7����������'�
������dK�hY�@���rq=����xU�Ω�w����:s�=:U�}��;'X�>r?1�fG��(�9lT��`����'���w�`��s2���<��5����:��~`�D��5O��=��N��*Ճ5S|��h�\�����dvǳ�S
*K�d����d�N�����V�84�w���@K.�j��v��%��g=I���Iw�]�T��hqaZ�&���V�~j��l���ׂ2�х��g8�ױ ^��b��TxW{iVC ��&Xw�N����?���#�%��gzɏL�����ۚ�a*���] ���A���Π�!���a6DJ9^I��m.��s�H��FQ�/��\`1�Aq:��*��R�,PTq�MМ�:x^ ��σ��d�M����K��k����*����)��	=�'����g�[1k��Lˑ��_+��V$ZУ�wj���'9�.Hwl�#9$�KM�¤O(�Ig�e0ݷ`C8�MX���vc�ؑ{�rI�B �������ʙH/�����'���KXC?�h��j¶ R�dT�T!��Դ�0/���C �'���G���8�A��<o�~��.q��}q[!���~@L��eR��H�C��T����Bg�˜�C0����Jص  ������\� ��I(��T���˿�������5�J�ݫ�Y]��ĉ����G��y_.ׄ�,M(s�{������*��S�:r�9l�+�1��,Ln��! �8���K*d�!%f�	�c�u7�eP3�Ŕ&Z����s�ЌJO���:�~F�vׅ{ �� ��e�h�a����(��u��4*�zE���dSNV���{����ѕ�ܴi��h1�����0�!P���}Ǿ�lDx�A�+��Ϝ�����)���515i˾U������W�b�G����bw4���I��H{~y�����/���???��ߝ;G�4
[��~/+�{
<~�M'�����7�ףC,M��sX��mjgiل5=��e[�$��!	@�]��Agpk�p&��s^��o;ҫ���0��'��ke�V4��Ȧt����(�S��.ܾ+�����x=٢J�h��Q��G��ӱ�)"�"���+
+F+{��@͸T�1�%UU��j�ێF)�Bumoٍ�O_9��5���Y�$�B���c�-0!��8��eL�z<����n��F]?jm42�]E@�9��Zn�R�ѯ�k@��O��O��eʌ��Z��'t� [�)��k���~���p��*�;����쭓��/c�j��^ʣ�MQ@�TS������.}rl��� � ���{�86�����[+x�g����!<6�ˬ����؛��B�;�#��r&���yՊ%x���>�W�Ǒ*�E��9���ӌκ �_�Y�۸4X���߿��@�e�^�d|>Ͼ�㳡����G�ؖGP� h�h��"�ä9Ջ�"`���q���\���Gr˦^�
�~�c�C���Q�`�>�)�?M���D��T�+� A�N�YU'jY��d�_�_�dӍ�H�k��I�b��r)�u^���� ��`Dnq{���=jNU�e��)u?hDDU�a�gutD�VS\�s����6�$�zgR�)�-VǾ���@�"���Zo��$0�4?�6�on�[k-y�R������y_�VFJ�nw�[�|�(��Et��>�"k�g�i���H Xotp�Z3kx����[�MP�`g�K*�J0�Y "J��5ª��0�-rE����q�1b�(f<�;����߫�^+b�QX�I��W����s�B����AJ&RΧ�y!6����;�r�����%|�s��6�6�7VK�f:�$�@�K��f|W�z�O��rqK��Y�>��/������
��tGe���-t	1��}��,`i8�1�f+�#�f�{�֬�bu�M\��fM���# {��8����Ș��QE�A���e���"a����s�3�F�[�B|z$q#��S��p�����x�]�= 3L�����D�QA��Kd�*Qw�(�f���:>�*!����p(�i�Zv'_��w>EX��6h�D�Y�����1�;��a^�Vٗq,��#]���f�xd+����V���:��Ǔ�A�I�=	���2jBD��ZaC��[7�M��%,+��� ��G&O�3�M�?N���=������r��"������U��"�q\�`�.ڦ�h��a�R'����g�~�)QA��LV��Zթڶ�w�\�.�#0Гq6h<�O�  �{�) "Q��gJ&(�Ղ�Jji�uCFqH	�j�Hz��1Y�ʤ��&����~�Π$01VN��gQM�="Ъf���cz�Z��#F�=�/��? �J��EzI�6 �&n���¦�WB���"�������y?� ��#�����;#hKڹ��7�a5�`���ڗZ�w+d��iC'���V���8~'W�9�B�C���&�u�3�/A���*�XD����Et��V~�:4"v
S^v8��.�[�JH�2�,_����#�%3]��6و�9�u��Ϩ�E}~g�}6"��~�)r�5@o4�x�ꒆ���t�>��_�f��wi���߬��U%������?�GB�&r��N�O��<�@~��*�!+G$Y�-��J�6���ԓ!���^�E�ЈN�h#Dn�O\�uN}t�������>Q}�
�fu4!��EV=*�}B8 �⋺�����,^�d�_��	
 P�a�r��HV�-E?�1)�!~�uQ���
��S9e�=@���9�t�p���g���X��i�
������6^c����nn���a¼{0W��sG�&�<5�Ə�s�,�v��� A�������l��]���mA��EA|y`xV��U_P��f��`?�X�u��/�7n��Z�j;n˽,�Ktz ZBQu�]��ƨ,�����}��D=p-{�Q
k�t��A�4g\BΜ,|���v�`�V*`�N|�=���[�B���(�R_��_�uۅS�UKe��Jw��.�,H�;A�
�/�o��湈\b"���% ���#���B<^�B׋�Z��j*d��O�w|h�ڣ%�.�r�̻.MB���6ף�B�:�,b�~���HR눤�׫����+Eր�=mN�x��@�;�c}�����V�Q��y�Z��y�+���X����I���]X�+��J/�^�#h�c�܃����8�ō��?������D������.I<Ȁ��~PAM�&l:���Ł��1��ptH��b{�F]��&��u3/'�0h���Z>�]7��.�vbӔh���`h���г��A������ܾ�g#�%��Q�Q��/��z�*M�Ŋ��p�ɀ���k+:%$�����/rxe��_�㿉Y����?p��t�W�"G�Js�"I�F!qW8Q�#�
�*�,�s��N��D���~�=y��f���-J	f�e�{rH�P���>�V ���$��b�vZ7�	NT�g�0xI=uP����<O�h�:�^���d�(.aŬ��RƯ`�2
������6c��g��"��T˻O�@	)�j���~���=f�&���IK��k�@�O!�j�����aG}35�Y:��S���x4�i�����2��S?A��<��t4rfL�m�x0^6>]u�:�;���U�i-�C:���H� ߭�LC��GBA�(7�N{rm�d;�,���,h������>Ӱ/�?��6��q�bzXN �i�r��d\�"�����( T�	�A K-��J�Q��{�3wq��RI�������i���>Ħ~�D�/9�/�42/%�S��%���$��n�2$����u%��n���r�>�}��H�����.��mq�j���?���zK��_�M]����S#�9�s}�4��zJ�P(�:5�0��DG��H�r�q5�UH��i���j?�Yke��t�C!#�Z����΁�G���k�CD�&�r�u֝�+�h����So49*RA��p���S��Y�%��ilx�'��51����ї3[�V���p�0� �S�k��#�Y�Q-�����&��.t[�����|D⻃�j0��c���Y�(�%ؽʸ2M>U�a�|��̬kFл��ݭ��<�kD �����,iq?wf~	����p^p��<H������a�IqcG2h�w��y�&i��j-���c?o��뜸]���]�6���X�H�@��24Eݮ�+C�-��6cN@��Y�����*�-%���rz#����X�X������;��F@��HbRT� �W�"Z�̹�H3J#B{�{�B�L�t���p��i�p����k�W��'�
6ѡ��YR/��4X
�ʲ*��1׹��.	ux*灙^*�z�.����o�<4�G��8��\�瓑ē��OE������r���:��B�a��&���
$�s��ܛ��,%��T�΢�F��1ӽ����yb*ǳ�2�m�|�Sۼu5�ʿ�="L'ח�\����Z���FJ��fU��k�]����L���o�ک�}�A�"!a5�}�#�v��g�?�;5f�q���&�<}$��z�b�������7���.3���ڜpQ.��1h��r#6b��S�I�Dοa��(S9n:�bl4��[�6����T%2NX���V��e�@-jo(� �Sl��(��E�,�Z��H����8G�/_<�� r�.�ݜ�[0�
`��N>��>�g��$o֊���37p��Y��q��6�����v��ן�o��{�o�Ͷۺ�*R����ǟ�s��:��(|ѕ��9���Nw������M�ŉ�kX���	Q���c��|PiZ��YI�J�I������-�dw���Q�g"h2�h�,EJ���w�O���x\#���3"'Z��Mm0�����46J��\�WEq �����ݵ�X)ƨ0N�[����U��@�c4�"C�)��^aƩ�5J�+�2!�G���Բ��9h\��ruM+��Z�3[�{�`�R"� ;�'��4�b��~dn���:���B�	���#���"�u6��1E�rG�(G�G7Gn�w����:�T[_�5���(��g��u��Y��M����G�W���zm�����_E�1$�w��-�]a���L##6R�/���Tes�=S�B�i�Y���MG��¡L�>M#�~p���^��O3��nz�
�MS9+���@��D��O�Dl�������5�Ϗ4ά�,d�gG	-��&7�����8���m����՚�d�uA9� g�
�|U���DXq�V��_���^D�/X$kQ#�u��Z��:�\W�*�	e#���&['h�������A7tۂ�:�GI����Thq�B��yU���`,m�M�̓�@���*9w�aMl|�;��ͯ��	�Q�NǇqU�9�D��Qqj�*���B�b�m�*H�ͷhM��>q��ŽF8� �u�x�k�k����tF�̢c�ĺ�H��s
���_��~o�)Hҫ�s2D�D�a S�����NІ�$1��QM�գ���)�'����ĺ�Q�[J/��~v��rZ���w������=)w��e��+��cnBQ�\��}n[��L����S��r���ֻ����T��,��c0}�"�۩@����31@��_5�0b���|��K|u����9�gMwŶ��Z���g�@L{�P�� onʁ�%��5/�o/Y1|5�	��_�/!����BW�>PT��������w& ���4�l�Yj�ݗ���1Lɀ�[@����"C��ܥX�(Eq����&&)�$L�Z6��JP�/��&�����tע<�٥�Sk�>ie��3�ĳ���o@�W�FG�j~���/���
T,�s�lE�<��i��q�� ��- xa���ߕR+?�C1�b�IhH�R���u�(��C�
y�W��u��}e[�*h;jA��ˆ�~@��T�w����{�1�:��aB�g,+p\䠞�wo,�.���X&����Eo�l�wTι�Vq�q��D1�GU�,���/���fINj�d�`��}��TK��"�s��R�/��f����Gv���ˮM����h�Q�r�X���SHQ!F����T?������ƭ� �(8=̔��
x����
㯳��5ұh���ٵ�<�sD���?��j��aO!�2h� Z7H��Y*$!�>p�󜃒;�쥽���3�3GB	jo�Q��Mq��D������.)��u�`������=9�݄T��ۿ�0W�w��F�����-Da.5xEm�u,��
��1��n��R(��T�����cld��D.�A�.���U�^��m��8ٿ�c�V\?��qD`�.w$��ݛ�>�퀑T��؈�y&"�A���i"5�s=Zٜ�J7���(z]/�����o2f�Z�`�`�O� 
��@�p�6�������N�C���BFQ��#���`'�1!�#��8��{=Y��YG!ւv^_��p����ZQ����q��!P[(��)�a-X��n�~��ȵz������!�9q��e���΅t���T�0�#!P��C��)�y��Kk̎�B"7-�ܳ0�)�]��͡mn�9X-��Dn,l�R�	��D�?���uYv��̍�����8��>�����q�s���F����ђ�|��O�ٗ�{���mrW��]\c
lD"�2��qt���/�ӈ{w4Q�{J*���\ �_��bŊ�o��T �K4�Ԧۙf���I1�6ua�K�;N��ɽ�E�]�T��~p}��x_�\��ɴ� ��_���2+�HK�Ŀ�֗�}���& ��p�Y(§杵��l[�v ��� {dKy�{�e�$A�����ɕ�~ՠ?�i����ed�qp�X_�8�L����v�����q� l=�FY�^���zyU}X�p��G�&C�b(Y�,��!�x(rX�(Zq�#gW�6��Xը)?Գq��"�C�h���'��"�tL "pyƄ~0;��6X����Qk�"�S�#\5RS��:�5Q,�U����?���z�������b�~�Cy�3��I�0D�WF�(-ڕS�#U���a��<����f��+Z�=�"e��J%�㈲��~߄B4�۵C�������~C�`��~m�8�?��Yܷ��t��[���Zu���17C��f���ѸlI{p�[�J����[�=��ؑ�o`�PS�>%{�|��K"��̜�-o����G�VU���$�.4S���:��1��s "��*D�"B�7��Y���ec�U�܈��f�7T�bm���a��;v��?��\�Q��솰dT�&"I���@У:��>A9�6X~ͽ�X
���ǝ�WG�"+a�H���N��i�@�Xn���mn�b�bfr���z��\�L�����1�#�� ڳJ`Q@�M)DO�n��W�OW�n�v�+�'�1^�LX���UV��w$��oXsD��꫍�^d��9�������=�sQ"j�_����BD��

p' ������x�d���hoڣ2�]K�{�5x0�@,������J��T��"�J�Z����u�~�w�3$B�{k�b/r��G��q����qS,�4�������<�������_B�+���0e|������/7l�x&ꑅuI.w���C�7ø])�:�p�2:x�ѿ�hi ���Y��[���ў��5Y}���_Nͬ�5n4�wR�_��gև0�U���: {���?ʓ��|w��������F`�T���A�ʄ.��̈́Z�J���Җ���)
ѵwI�(et�Њ���Pa��2=p����C@���|n�ظ���o\�V�.H/c��y�|�vP�D��w �}��G����L�S-��Ec�0���WI��5o��n������n�[��������[�Q�=?-�$�/�ˏ4!��k~�-����Ί��8����X�D$���;@%���m{w���OT]ਛ�*� ��]5F���*~��Wv]�06�R�q?W�W�p=Q���9ks*l�s:W�<H
��\Cg^���w��lPˌ���;Œl�a���(Yx��H8����CJ�J5��'��6g�N4E��$���\�0ո�������#��q��~4�Č���޹�����������eC��Ԇ_�Y�Jl�#�4��X�^6�&�˲���Q*٭�?�sam-����}B㮶�L`�����e.Zn�A�� �&-ψ�)��I��A����fJ��qOl澕2��	ձ���ޮ}���H�ܽ�2���.�U� W1Q!��:|���K�3ƽ�.]���Lbݏ���R6����n�~D	Q7ҒU�w��c�>�sCS�i����AL��W;�M�R�g�����!Y���6e�fZ>�MlF/�:S���RCWl���h�F$�y�*��zZ!���?���Kt�J�ߎ��>��c8�;��
_���p���;��m��6dK����q�U���Ra���8CvV }���b�4�u�����%��@�	���|�}LP�]�X��I� O�&�#��*�ԉ��*g�=�L�B$�$:�΍��4#d�����z��M/9F��Ȼ�^��m6��㻻-�NG�(%�Q �xVorjI���SM5������
=at6�YƱ�d�h�h����{��n3ʨ�8#�� �]��r������*�� k&v,�h%��
H�9���[3<�^Q��eM����8UŁC��m��ƍM��#�����ۻv�#m����+����Cznd&�m��]��x���f�L���P�Hj��QL#�{݅����������0~H�����4*{�G�����I��m yE��	oq�2�������ﳃYH�)dˈ�e\6�rq=�P_�s��r���l���V��Mv��3!ͭ�N���x�Jѓ��h����o��CKiP�:!�x'�h�_��qhO��IT.�� �%V'SA�&$y�˗�;Q j{A��a����9Q���c'�[�P��c�v�������z?��u�b}����ް-����uJ�7t��1����pF��/a���v�C�S4�Sm�r]A�1�p�����z.���%���{cC�++��(�M�o�@5�;�Y�1�A���E�����q�Q�>�uv�_�����|1"Z�b���~o;��z{�Ḳ�A*���T�N#��L����%�v���Kz����\�����כ���£/M+��up?��cz��:���e�/�aT�hz�n�7��8`���E^y΍-��/���V𐏲��׻�,��4z��Z��ɩ��%�:h9&�����a�>�/oeV��?�a����D��0C\'jZ��D?S��n|�Toe�X7�����КWF��6I&����U�_�V1��]uD���j�n�`�R�L�;P�m�|<��Lp]ݤ�%2ZH}��1h��9����EP@dw	YJ�>m;��E-���X6a�r&[��j57�c�4�_\�+�Nz��$��D����C�N�i�SBg�9��H��he��\��8��2��aɗ�t&��>i}ʘ����Q��0) �e�L�OP ���E�f�m�2�0��Q�~*��b�;�����ZlD�p�����j��r�@�>z�O���8n�gq��.q��8�?��7����A�v�����95֋��fW�/�&��~?a���^��I�@U��
@�h1��(��zڤ��􅼁��{�A��iI����攎I�4�v}���V.CX�b�@;:@F4��*Pq�\�����W���sOgB_���j��8ܨD��9�|��V�wT�� #��H�= ��B#y�qW�q�W:�X 8�{j�o�\��ۉ�v��	4.R�}�"= ����(1)�ٔ��J���������_��/U
%+(�篆�tJ?�ss�o	S�z���S�d��C,��C*[�eV�x}+g�QK��{�v�'�Qj|�ѿK�(ցF}�g>��f��j%���Q<����[tA5�Z�yq�2��v�n@6�SDXi8��A�ͻ|�2<a�:�7�~�X��n�J�݈���p���O|��9�w���P�jl�*˗��;�bl�$@>�g� sߓ�6��e,�g����>TA�`Õ�A��x�e�e=`o�]���(	$΋��( �t@�Ql�|WA;�D��N���l¥�L6�QS�Y�s�վ��aP��D.a��)�ˮT��ZN ��nG�y7�>׃����f��r�5R�Z�Pi��S��6z8�����,r��SZ��i�����15|��+�_�{����w)[IIP�\&BT��l�$ш�e9y�o��R*�l
�G��E�[&.;	z�2��V�$���owp"iZy�^\��	�0Gڞ�
m3���˿���!>����������o�����|}�?�����������o���~��������O�W|��W�����=�������������~�/��������5HNs�& 