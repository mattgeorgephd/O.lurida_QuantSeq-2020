�      ��	��GQ�_�{��sf�sf&�$���d#�!g&�00�*�,�a�%���%�,	
���� ��"����u��ʅ+�^�{������}��>�����Jo���U���ݗ_��#��="&�����B����_���|�=�y/x��o�K�߳^�§=���y�]nxa���}�dX:Q8Nd>lpI����Di�
���=����{���[L`���w/�~����ي�g$�ގ��!}ҷ"�����4��|�&c��~;����)���d���o�[��f��o=*��t�㣥ȧ��$�'b8~wL��Q~���5~������]�9=����}��	�xp���`�����^~wO�%>���g��	��o7���M�~[P�.�O��xl����B��L�����*ܜ����	�����G�'�܇����V��M���CzH|��;����b�'Y�d��\���൸M�����n�������_6���w��1�&�@�Ӑ__���_�7D��u��iI{���>}~�Xl7Xm���}<4��������t��w	���)���ߊ���'�;�����g���Z�>?s~�E{g�^h���[��������︭������o�__�����P^������ϖ�����������-��F�l�[����i��m�?���J�?�VG���륅~�`��C��g�������&�w���.�k��`���	�����מ'����(������#��o��j�gK?�~'?g��}���t�������Z��N�G��d��1\?�ٟ�|����	�>y���^Г�M��;-|���?�:=�P����}���"�ﮤ<�)���Mҧf�G���>?�޼�R���$�� �
�ی��/���'��葭�k��{f�R~P��{}���K�����rR_T���F��y��Ox!r�����s�. }%��?6���E������4VOA~�+[?�d��"=�o����F7�x�v�|W��1�N9}��Ӗ��|�zwgR���_Ϳ�$������ϵ	�4���q�Ծ�S����������O���Mȟ�����������1O�7��դ=�����Y}j�=��_����#���{�����}����=��� L�����~������~I��?��gn �@y���w�w���]�<=�������[���{R?O�/�(��[����������ǫzQ��A��ߗ�^�z��uo0X�����뉖?��U_f��-�'��%�㻩���'��>x3���xz��a�z��ۣ?�Z�!��]~�^/��o��@O�ߧK�n/,E�?���{�,�~�$��[ڻ����@~����?��Z0�높�~1>~lo������7�@^uKI���K8_��?_֯��i�o�2j��_Ϳ?}\�K��!)߲ǉ����q����$?��Z�C���p�z��+��'�w����?9�j��K���{�����d��<iO���/�k����5���ޑ����}	��~]�On��������=����1��f�V���d:a���{hﹿ��П��y8�/<���N��ǋ���_���zV���:�oo�����7"_߬��sAO�/�:����oK?i��_(�(O��O�1�?҇��<���>}�����/�|P_�$�Q,F>����ǽz��ׯ�����1ۗ,���]Kߊ�3�`��������-)_�W���5�u}�Е���O�~���]_����s�K>8�h���v����O>}}��'ў�z�5��_H/����y��U��!��-�x�����x2��=�z�^�ίZ��4�ۓ��LB/���[��,y�x�/:=�Y���L�;E{(ÿf���n�_�??N�T�>�x��R�����q�e+]��^�_%|?[i.��W>N�k���a<�������??�v�Q��F}\��>o�Ve�d�ޯ�d�t_M��x��Z�	�=)%��#ڸ�^� .4�v�>�O������-yN�x�Ƙ�a��s�X�3Q���Έ����g�yC�������G��NGz��2b��Q����	��gD㛝~��^c�.�_��~���xt������^�WZ��C�w>��^�2}���Q�����~�>�?U>��p?��W��M��|?��)�2z3�\kÓ���������/ߕ�����H`��l�\�'P�R�g�G����46o%~�y+ߕ��&�%?��P��ΏZ�y�����GD����z����C}�(�_m�(����ݧ��Ͽ������b}��2~E������zi���k���g����&��q��8��z���`�����y��<u}Z����G�|>��ؓ����6���uzH�?�`�o�e��^������k{y���]��H�����|,��s�+~}��E?��#"��.�r�H��W�O
om{?�g����p��_��gm~ܜ�Ks�\����%OJ�Y�Ȫ���oj����/�_��S,�s���r{K���?)m����j��/i��0�[����KzR^i�~
���������ԧ�k���u��=��<���U�?*���O[�t��?���߃�~~B�Z�|�v��[��{#�7l_�;���W���?��ć��Z�5H_2���|s��y��x������c����?0l�#3�ض�g���鷫|%�$�����j�^m>���G��V~Y|�b���l�xz�? ��������xŧ2�!��[c��,]��_�/��<�����}/O�����Ӥ�'"��5�F$��UP��s_�Onߴ�<�Qh�}�m�W2�������)�=ɿ���K���_���7�o�?�����.��}�g���[ryY���$]����od���_���z�o��>��x�_p����N�i�3��j�wXu�?@��N����|6��_��e���}���_��e���>���~YwE�*^g<�ק��'2�K�9���������{<�����|P����u����zS�_�����'1�9��o4����'ɾ�G��Ŀ��}�f�#�N/�u���7��wE�\�h>�z[�����(M>"��&O�/lp�/|[a)��%�����~�sR�b���.�����O@��}E|�����xB?�+��/;������1��e��Y<�5���ȟ��/�o�������'p=��k��/�k�jo�:��E}���G��cx~��G3z���p=��3{��R�����l�Y��<���_}}2�����7&�����?��ފt������G_��Cu��"����#���ݷ��g҇�u1<_��[�e��!���y_�ۯ�������[�|�7W���WE��?K���u.F������j�����K�7��7�}}?��E��9��R��_��;�>��6G����h�����]��ףO?��C��G�5�OK~���߅I~�����a	�m����'9��x��> >�o(&ǯ!=��_'�G��e�P���do3�����>�s~8�3���79	�zRӹ>��'|�󆬟����˳����7����gy��Ke�^�x3X���}�6~������_e]���EO�W�v���\�3�y1��>�K��s1�OD��P��<�غ���K�	��i�������\����?r?��Ѿc��{cx���{�?�fR����k�{f�l�����l��=�|nN��o��Z�cC�0������ퟫ|��$�j��k�#z>W����8�����ύq|5��S	��.?5���`))��BR���}�H��������/�$�~�~�?��[ +��3X���_x���O�K�v��x��/j�52�i���i�����f�s�:��O����F�h��9�����㱝���P�[t~�D�?���ϳ��O��C���N���Ǿ�'��[����ۖ���Z���`����>�{N�Kn��{��E���l1��,Y�����%�{m�ǚ=����G:����Z���w�����B:�)o��>�ٟ�__�'no����Ͻ�N���7�W3zJ>�|-&������������U"��͎�O���i�;�3f�u�����飾_����(�d�1�io����{�8>���hoJ����_+2&8��P������J���y?-�l��-}��CX��}����W�>���K&��������#Y��9�j�^�iH��F��O��];���#{?��j���鮟��I~��{���$@�ˁ�>���[ɛ�f|��ߵ���|���"@y���[#�OF�^^���op͞YMꫵ�ݷ@~o�}R{���:�s>	�3c���<f�9�[��\Ľ��e�W��b����_�W�O~+���뗈��uz��W�ӽ�����:��/��{�����{[B��M�ȯ��/��c�ch�f��J}������x����?�_�u���.������sɊ�пL?��4Ɵ���x��O����6���⯖c((O�H�f<�ʟ��_dEwf���k�S�&�y�!��������y�e�/ޡ?������}ğ���3�����d������{M��RBO֯g�X��3Hw@����GN?�/���_���M��;�~�~�&����Hȏ���!ӷ���a�+�[��h��^��������5����?�j�����>9}W��h�K61���3���A�Ivz~�$?6�g{��xP�g�q�_�ߙ=���蠯ֺ�7�O�h������?p=V��� &�..��I���G��ɚ_�7���a����x�/X�x��a����@�hO��_��k���K\�:�|Q�Y|Ö�7���W�א�N������`��Z��$��]����$�Ӟ�>���%+�����-�����/�?��]��~j�M����+��x�Gv���?n�����eIz�L��{O���Q^�/W�Ѥ������%�k���K�:�w��d�,��}G��_��,>M��~8P����?\~����?
��ⅉ�p��S�4]����4��O�����ث��Ex_�ǣ���ˬ���t����$}#曟�gf��/b�Y?�� LZ��ϙ�����k�_��>�@}^����I�����_Y<4�+��o�C�_ܒW�F�����Z���K��Z�o�S�e���@�!��Ai�/���,�6��s�_�>?��p���ۺϹF/K�+Ɍ��|������"���}&�����|�xG�s����xo��4�����_z�~o_�^���?�������%���<A�=�a<������3P>;�E����������á?骤�Z�SԷd���~I� ~��9�/�/�e����K-}6��w����߿����<��������w`���w6�-1�������If?���_2���3�_u�l~/V���Y_m�����h�Rd��B��y߈�s���1�������3-{��Y��~���O���1~Q���F�콣y��Z�6�ϟ�������O�x�~w�,���5��o���k��p?�~>����͖������>���^З����,]����
����{ٴo}��~�OE��G�V��_�?o������U����e��n0�sa������i�+��^����~������Z;�Gu=0Io�C�����/~�� ��y:�iB���B��L~���x��Iy�g����?3�Xu��i�9=+zCR�B�������~qy*���.[���[�����\|OB�O׿�5�����?���}����<�e8��,_�y�g�Ou9?�>9�?�o>�Tq����^���K�߼ߕ�\˾o���ȟ�s��#yy}}�"z���P�0�=��p�ǥȟ�ߵ������g5��P�!���2�EK�;�|y�YM�y:��z��(ߺ��i�1^􎀳����L�ܽ%I�v�߃�yމ��������v���-]�9���|}6k�"�\~�z���C�f�ym?�����;*���t��c��M1��Y|��K~�c˿_[OҟA���G�����xW�g���,O&��
��� �l�d��z]?�_��e}_�?�϶��p+~���f��OG����Ƈ��xww+*��ȟ�7�ܷ��`s�� �{#}��aj�(���}Y�7�?�nr�b��P�8��T����3\g��^��>�v�{bh�e��@��V���� ?O�n��KŤ��*j���߈�}��y��>?h�=4����3�W�����#�O��ek��%�<��~�����C�s�Fy�3�G��8{��F?�����4v����A�y`����!����zS>;}ն�����_I�R�������Mk��>�����餇`�ǜg=,y�����,����7t��Z��z~i�*�OyH������`���Ճ���ǳ��+�ߥ|���4Io������c=�?����g���}�����_�{�1k_?�(��׈��"�/�~|�����[}x�1�?a���d�?�|���f�����|�h����j�O}���<�K�} ����P��^2��ʇ������W�{7���_�����ˋ�������㻤oݟS���o}�$���}�o��x������I������r{���<F�ҟ��w-���W����R��<n6��Պg�������e�$~�䋀O��9I��3�g���G���G����:�w��C�>��X����%]���5?<�D����W���t���?�d��8�����H`��'$�o�"�%�0��ij����"�=��~v�9�;_(k�3�5��~'>�|��Yp&��!�����Vޞ֚A�>�v�P�e�gh���۞�����G��>\�������:�C�ǳr�6��%���	�Q!Q������ ���c���Os�X�����X��ϯ�o�t��"~3�uw�B�Ko���]��]����ܣ�������W+����~��<�|+���ӡ<������?�.{�ğ�|Q~�0�W��[���&���kv^a����;���8���?Q�,~<�����"��%��7�@c��,o��������!i�e�)L"�?-�"�����������~����k���O8������x�}i��^n�W��߲���=�Ny��f�����i��������9�������R�Ǻ�����Ǣ���5�yT�����ez����￰?�/�_�����M�'����k��Z�f�������UnH�S�|�����}1���x�ho������?5��F�}1��p�6����ͣ���~�z �G����\/��i�[e}�����$M�����Ki�{y�C�KD{������g�Fn�߲�3��޾�_��������1|�:���~�g�q-��e�/�.򡣽�����7l�R����-��Z����=���/v��d����V�g�5Ƀ�!��C$�j��^?����h�p������g�x�?�Mx�?�5[P������ӝ�$����j��C��#�ߚ=�
�y�zD.j����K&k��g�g�e���b�쏯W�_\R�|���ۣ��0A��}./%+���+_����L�ooF�l�Z����/�����N���.���#������0��}P�ov��	)��|x���/���X�	�C�3~Q\��V��#��m����<鬍�#��'Z2������3}��Hw��"_�k|.D�����ݓ|����7��k����sIy���O�X>oM�?�{����,��O�O�_��"}�sN�l���ڧ���1�� ����d냒��?�-��`ɫ�(?�����	���i��À����~(s��鎏��kAσ	�k����|��Q�Of�r=+Z\���~h��N��A�?Zpk}�)��������0����o/�?J�t�����ik���/��؈<3|�[�N,O{��˼�y�0�oc��1�c�޵x�,�������!��z?1�/�3j�3~4����:����Z|���P�|@�~���#��p|j�q�߻��~�x^Fug��1</�� �~�o��L|��f|,�C�O~g|�w����r�J�:�Ϥ<Y>�Wm�9��Vw��x�7�x#���aR��o��63��������|��d�'\ß�������x� ���d�?y�
��/S��ҧ�)k�vxW���1 ��1��y~�塚|�-�Ocy����������,�V@��������ޭx4�7���y\�?_����<_Fy��)�3�G>��/���7߆�f���|?G�~U�G�>5}�p�����5ޯK�������\dO��h��z��	�f4��3�ǥ�%}O���Ѣ�J�=����_e<����E���W_�Cy�EwO�%���'�����P�g��|�>~�_D�(���j��I~�z8,�����稏��?�j(_<]�W&�Yn�7�/�4��=2�^��^֗�1��jl���X�w��C�GP[O�̞#}6�o���w��|^�y]s+�Ϧ����S#��S���i�~��s����|�틿ޅ�2��4��d����Fz�>?��`���l_�ӯ&����F�#�?�%����U���J/O����)��������˒��o���b�M����R��{�p�������������ޗ���������H��׊�Y��\]��`���߼� �������$����,?a������s?�lN����c�Z}-���W��t���Ԝ>�o��'�Wݥ��K�oj�Ŷ��$��F>~�_��o�Ez�������	�y��^��_�'���S�zwԟ��Z�c��w��|0���X="��ۊ���$鬏�-��oK�雯�͜����l�Os�����O5z{y�u����o�Gԯ�һ%����vW������G����߭��G�/����D=�-��l�I�+�%����d�By�ҟ5}O�K��&�H�f�ى�����>�7��^{����㫳	0�v?���������d�O{�믖<'����K:Ə:>{"?O��[�}'���yL��]��c�����CT��G�~�֤<�O ?N>^I��d�A�[�91�O���f��~Ώl}��?b(�Z��^���ػO��I��}���#����/[��s���f������>��U�R�Q^p��PҞ�O����@u������?ϯ��x����g�V|3�OD�������/��gW�'�o���;�?���?Z~���)�}����pߛ�_�w?���O��������YB�U�kｳ|K�:LJC{���~���bx�{OR^��y_��o�Q�����ǟ���������Y���򴏕��;���g�����_��sf$�ǻ��;�oj}���\���Ӻ��=[io�z��_���ў���W��I~����ӥ����!���}���U�ϭЗ����w&�	?(��er<.Fz+�Bs���a<@����׼?�����o��i^{��ɟ��<�x0Ɠ�꟠��C~Y�gz��}X{���l<#��;��>��R��E~����-�X��5�l�<�\��-���J��w��5�G+^�E��Y~���C�p~�=�����b���'�j�9g���>�ݓ"��ÒG�{%��L^^���_���t�O�X_�����g��^k��_���g�]�{��_==?���.�����'ǃ��}{�����~�o�)��j�a���>��>��G�^�t�q�g��r�%b�^�����C�[���~Z���"r�������{j�+�������L�8���O�O��(��3���-{������X�=�S_��<�}/���l=ժo^yO�B��;�I}�=�?�א�ݷ��p�'j��.�O�b���c���l}5ksL�i���$]���)�?�H��y�~�������>����>���^�<�x���'$�%m�߇J�����W��٨�司:�����e�7��O�?�gh���!�:�WA���5?����IΌ���n3X��B�w���^�ɏ5��<����R��������w'?���~�￐^|e��m��/�S�?�>�� �_�����������5���x��=��ܽP~�����E��w�q|X�������̤>����P��Z�a�Odƛ^>�/�՞���{��jų�Ǔ�_xma��Y��ō	=�^m|��w���~���7�S-�#����`Ż^���?�������x���R�V�e_<2ɿ z�}�Y�3�ͼ�?�˖��a~���+ח�?�[���wړď��5����/ޏY�7���	勤O�t`��'����pw����X~��c����i�g�X�p}��Oi<?MzS~d�|b����k�;�猟����I���)}�����b��>��?���򮿧1|�2�����77�N�?��+�s�W��G�^�ֻ�K��+�q�`��u�';_B�U������~M����I����y������!���R�����r��Y���k���'g<�F�����w�"���z�Ӎ�}��Ώ8\�7[��I���Dˌ�6��0�}����k8���3�F�U��d��Z��?��������G�f�8�n��~�����j�g���b����>��\O��k��h��|��K7��M��|䧾���E����h�1���~�t��>�?�פ���Io��*��J��G�-�V}�Ogc���W���דt��߳}ޟђG�*$����n#�̟.[���zҞ��s�?���W��4�O�������(����Z�6�;��L_�/�_zH�O���G}���n�v�������G!������-~c}�}-��g�#���qz���<�i��I����(�k�������Y�g�tY�N��֚���e�����V�<������ʇ�1�O�ݯM�d	��>�3\�n����3������j���x|��1��vz���O�B�I�⣈/�\���?�/c�{Q_6�y�Cs�"��D��%�.���!��G��c���WО"�I�]߯c|��zҭ������5���גς3~g|㹕6M譹���o����#҉��o�~���J��IY<��2}�4??Y�G_�7��6^�_q�SP_�����n�f+~�a���@��?�K��>_o�֟�Wv~�p^a�GG>^�yօF{�+�z�����{4\Oe��Y�� �����@�OL��;�����O��M�����i�}��(<���6o!��^+^��!�������?);O[�'�Gd~���'�,O�ފ�{|�O���l~�����̟�Z�����}d�g��0ħ�/�c�����G~���O>����9�~-����9��tsR�<�3�>��f<-�ú�qg��K1>��O?�o7F~�E��x���g�/��@�����~w�_���I�}�k�������g�|=/3��A���Y����y�2��x6�G�E��AM~r���)�o�?P?f�4�O��L�(��;�3俕��� ��r8�їl_�v���/��e=�y�Ⱦ�7�Yj竲��V�2�[Kj���7���+�{�d�e�oٟ�| ?��s�����'�=I�6��|����~��7��v������R޳������Ս�)��=я�7�>�k��O��?}3�l)����/���Ʌ���=>G�s�$?�+��D_!��}�����Ë�V���?χf뇥=����ݠOD.���'��u��ͣ�����O���k6ݯL�� ��>�/*�b���'�h����������g5������ȟ�W��˓�[0��%����瓔�d���{�>ޯ<A{����/ϣo����HO�*�m1�'^��͟,^�v������x�>vx��قI���45X��!�/���������/n��y��/�W�~�|���������O~����{}���/�7i��>�j��YI��}��7;?I����K�鮯����/�:�}1�OxO�o#=3��t�#�=�t�z����R[Ӥ�F�5Y~�}U��l�N~�l=;����鯹����~c�o����e�u�(O� k��/pX��D��Q�i�q���h�b<�ӣK�{�ߏd���T����������_�0����s{Bk����9C���7P�_�pv^H��K3�JpO�t�ߚ���w?Χ,}K�����{�o����ہ�4����y��5{���|vxw��w%����E|��%r��%�	���_N��'��������;@��[�o)�� �{Q��-������+��R���`��>�,�x}ҳ����g~>\s����g��3���|-�������m}���ߵI{;b([��x��<�Ǣ?~�'�����j0�3[�-G�ء���M�[���K�7���P��﮴����-�<|�~���w�?�?���$}"r)����~�g�Ob�O��mhO�}R�Ӈ�7��'\�Wu}%�챨��*��Ŗ�\������σi�x��1�ge�)��5~"=}}���}����ۭ�/�o����~�����+ʇ�
���z��؉?H����/��2G}�G������1>����{ch�Ѿp|���|f}����Ny���t�-���������s��Loɟ�ԟ�K����z���7}���\�1������3���K�bQ��^��/W�k���:�~�I5y��*;O��7�������Y+��#?�G�:���~���J�}�Wr��+����$�4��ŴƏ�׏��`�~җ�J��M��K���O�y���*N�^��]��)�2���k�?�@7"��?��������U_ _�o#����m���|��'q|&H��� �7y5��""�����?���������q�d0���w0�w.%�wV�
�9�����)ȿ9��3wȟ��^��3�?��[�>�_/��;��q����E�8\k��ۼot����]>����v�������kŻ0�����|q)��_�x��Ɵ����m������c��������k���O&O6G_މ��D���Y�4�,>�{z�W�<��4���0�g�r�`�ӜJ:������g��ɿ��l-^��ŏ�z`?�g$�ވ����}h�ӗ�9�|��3��y|9���~�V�D�?D{̿j�d��'��Ǆ'������ {��������]�����=��e�<�����m��i�3>��/��.��m�7'}[��/�?C�2���^��f�h{��?��Z��G�v~�{O|O�5_j�]1X����0^��o��;�z�!I:㭧1��%�Ώ�w��?�}��$����d�6�C3��ч�3�����k��H?��wE���Z��_$�	��S���J~f�>�w�$�5��	=�����
�o�$����F��OE{�?���I:a���q�R1������g��_���x�B���1���m7�����}�|k�'��?��R����a|�ӿůlO��k�*��[�w�g|��o�������n�W��M����v�ޜ���| �y�C��6~����E���F�����V��(�s��?�J>=�9�W�"�3�̭�����~���<�x=�ǝD>���� �'Cy����}.��{���G}��>ғ��^^� �a>~{���va��a�g<���>O ���{Z��J�ϻs=����D�L�ld�l�E��\��-�G���(���X�Zx�A<�H��������?8�j�Q���	�G���|����؞��;����P_+^,�?��W��<����/�
�?�������we�m�0��?���_�� o��'�����oi�_��:�_���m3^qyB��훝1�{�|f��+ʋ/A�<�����r�3���u�~5�2�Ҳ�X��器/����}<�>���#_��|�l��#�ϭ��k�e�giY}�?�s�o����3�+�>-z���λ����y�C���=ſ��`���˧7ʷ`����?��~���,��i��9�/�ǚ�7���[Q�9������g�<�K��3� ~<���\@}EN.O����P?�_���<�d�ǗNc�寮��N�����>�Wn�o��vk��I��K�g��xߧ���������»�r�0>��6�OFy�	<���?��?�T��s���-�6����/���Z�s�g�_㛽gG|y>N�d0�~>~��n2x��_Wx}��k"��JfϭE�~̚=���^���#b������=������O,k����g�\Io�Wy^��i��5��:�GV��2|6(��O�[\�x�Az�於����NݝK_�>��Kڣ>���÷�3����m1��F|���'��=�V��ԗ�ƣ���y�t^�}s����-�_K�k�1=��d<�F�������?��?���׿^@��Qs��i����O������K�w�x+�W���=9�Tv����ZR^�_��������Ͽ%��kN��������n��S��zC�}+����{��gE���/�1�����?^3�����>Jtj�>��_�l��xy{-�oJ�ٻ�z�v��a����^?�3��S�=�N��O��O7����7�G����<��~Q��i��� �N��~������}����{v��˖������]���w���\�������/��`�}}������� ��+c|<���r�B�s�;���!߃%}&�3{O�o5y��L�oiŋz{�v�W����u�^k}BX���od�������MyHy�᫺�~Fɪ����ϊ����^�%�Z��E���n_+���,���	}8^Z{]��V����D�G�?[?q޷�^�ww�q���硽޺o�aƃ����[k�ܡ|����aɚ�=eҟ�sw�����ɨ�u?�y1�����W�~~I���\��<���3�5}����������Ώ��3�Ӣ ����gh~��[�����/`�O��;�x{G�?�L��'x���q�k���[j��}���1ޛ�C�ֺ?�����y�������2��'c��{iA��.���3b�^�=��}�������Z|ׁ��}}zwE>,�t�e�!����^Z����?5Xu?��2;���ٚ?+K��|^����ZK�����_��A���39����C��������_-z�7ϯ���{�*���O��~�$����"}8M�od������W���Hy�|fI�g�G�����[���)�g��Y�5��]`��g����o����'�я�5Y�����p���-���#�L߈?���9%��#ϗ�����/Y��n�'�/,���V|z+>E��4Xo)|	���ٻ��x����L�+�O��_��W}m��p�nĻ��#?ӞZ~�ϝ&����3~��?+������}�{�/�/��3{V�l^��ߚ�п����/�7���xҿ��T�b�wo�����s����/�{Y�|$�3f���'��Ki�c&��0�s�+���B�K��!���3~������?�G�?���������~�k����	]��)��G}��"�.s�������2�/ڶ��5�ݿ������-���y��Ͼ~��p�-]��7;Lz�����r�Ɠc�Z�S�������{�zQ����C{����uz���g�����e�w^��wEzr��w���%�s�_1X���8~ķ����q�\���w~Q�����<Ul�������2uZ/=�7�֓�����ҷ�������}�$=�?�O��?����)`���,�٤~�m�ގh��t��ˁ���׷��{[����7b8�����C��������׶��{8�/��E�L����/����j��<����������p�B��x{k1_oO��xR���o�}}��~{���tv��Q{�>�B?��N�=H�|�ΧH���\����_�Px{�#�?R��G��YZ�l�.y����Ŀf�8���ߟ�c��k����hw�M��H��� L}0�!}��v��M1|o���d�����}�/���+hn�|���X�7&�i�����w��S����Gz���^?I�/��3��I?����}��x��`Ǘ�+�o��,~�����i��C��_se���;�[~��Hz��W�/����)Ǐ��?n����3~o�[���>�m�_S��^��~Y������{(�oNx-��MN���������`Ͽ���i0�~��H�*�G��D.I�1�r{���Y~^�t�MI���Z��C�1�ƃ�(�?�m��=��`p��.���ی�5���i�/�'ˋW����y�&��^���s�����<�����O{���\_G�˽?�?��q�Z�Z���'������|x��7�,?����������U��}m��~D~�Is�����/��M�^Y�߻��j���x�=io5����D��i��k���t~�l�:����O��xH����ޟ0��?;��E_�s��4��f�Ŀ��m�߇�?��^���/�d�$�'b��"��A6�ԟ'&�[��3A��z��g���?�_���8����,>�����w����^>�ioi<���?���];O��=;����+W}�Pd��sz���)�Kd����Qxy�G���>iF߈�{��7�������~V��N৺}?���������Т��3��f�վ�#�6_�),���?����}y����'<��g��_Ҋ?b��?��`|&��<O��*�7��a[��֏d0��4��l�K���}-��G�?&�o#��y�U�?VӿI<\��L�����V���oH��xG�#��\�Ky����O��?�nψ7��yyȟga������v}-�?j�~�������0ޔ��_���^q�&{�׿���߾F�#���{s�_���qzH6�<�������t�xV�?���<�F<�}ߴ%���eIy槾���{�=ޕ��g��m�����H���ӥ[ܿ4�c��c��W�I/�\)���~<����!�	��2����s��Q^�}O�C�k�?*Ig<۾
}�}�&�_t/)(�{��_���?Ƈ��x��?Z{����z�J����sP��W��7&�c�R���/`�7���s��:��������Ǜj�{UBړgG��i?rH���7b(O(o��d��Q>[�~	�����(ߩ�|�Z���w-}�U�a�d��j�v�gs����	����~��G���F_��=&e.n��C���~6���c��yy�*V�~�7�����O��#=j��f뗚|��;���"���W�G�_�/���qu6��h�u  g�w��g�||y_ǃ����+��|����~���s�/���xH�C߿��_�szR_D�y^wҥ;%���F�%�㝾ڻ���1����=�$�>�KE�ǻ��l}����?b��������2L�����:1��H����A�e�ik}���=���_g�|k���z{�{��_�o��*��I�ch�k����[��7����W���A��SQ��>E�twC����b�b����`��d��w0>H�����l}\������ߣ���f������y��ςu�~�@��Մ>�AO��ׅ<ܟ����;O�y�_D����U����<5X��w|�y��ӑ.��>�O}���<r��|�|8'ɯ���	k�^Oop�<�����g�����%?�kUx}�O��|]��yA���7Η�y!��$[����5��D���]���7���N��H���m�K-����!�=!)1��<�,�Xy��H�|v?:�[��|��g����om~@y�i���f����i_�~pz��d��p����H��3��K	g�0�ղ�6"_<}&c��������ti��	��m<�H��{Ub�߆��>��l����[���O���;��]>E����xD��E��	\�������ZB�0������y �߻��7��'}2�֚O���Z3�vw�t�k�R�g�i�K�?�{C��������[t�b�\?�>������ls��U���I~�����@?�k��Z��?���RK��u��.Џ�������x����p�o�����:˹p]��.��P����N�#1����P>:|e����5}��j.:?N��~�q�EO󧟘�_I裶~	����Ϡ��1^|/���p����jBO��c�yB�j�n��G�~Z��H���>`�<?�!��>��|[F}<1N�XlX���k��P_k|g}�t�rzӟS���"�gk<6�^d<���z��_��/����q�n��|�y��g�^^��ɨ��W-�8}d�_b��������)/��l�,��y��s<���� �U�������6�2���d}����꣨���_|?�����������>x���W�b~�����[������8�����p��C{�ۛF_����wl�Oz*��%�q���O�>���_M���X�}���K�>IK��ۺ�����o��i/{������x�y��:����o���K��'�2^����������������m�O�����?���On�������U��KR�6ޏ�����|U���|�_L�o��o�o�O���\�S?������Ol����1��w�P�5���Γ��~�N�Q]�h�G㓽_���gH����O�L�����?d�I��p=C|3~���~pzh,��{K~.E[^�_ғ������~R��G�_�������z@�����;�W��G����$��3��������}����>�����ׯ���O�u�#��2y��,W���S��F�6���v|vG>?h�о������i�[+��kO�[������?����{x;b��d��1���9���-���?�Կ#��3���oײǳ��Z�b6���d����=��>ڄ�[b�~����sCR���~}�ݳ�^f�D��ɗ#I�+ї_�M��~o���,�R�������	���G�o�G8��@ߝџď���?����g��(����I����}Ku��Q���%��Ĉߖ
�2�o�\^��#ȯ���������>���+���Z�i��oݿN���1���Q����|}C|V���s�~��_nO�=�_B����x��#�k�����֭�����M�o��;���I�<�O�ѿ+^�i����A�?}�wEN�k��?���+��s�G�ٗY<���-{��	�/��/.Y������xA�;��xط�8��WŃ<
���~E�u?i0�_�_�>��_��j��HO�g��`���>�Z��#��7�k�O���o��x�!���6��5h?�G�>�+�?0�v�
緧k�=Њ�yd�����ߖ�����Ӥ�y���k��5z}�Q��%�'��x���#�o�����殿���M�'}w����w$��W���[��e�'��^,_{_��%�=��f/��/���E�Y���=^^�v}G~���ϻD���L����h��]��kQ��p?��e˞�z.#�x��>���7���|ܾ��px)��?@���$?��݂��/�<���'Z����+�w���L�d��i���j�׏[ch/f�����5��`��}\~J���"�D�>���S��w�?Q����W�����+���xy�/�/3����}5<�H})�`�_5~j���5ӿ���[K�����w4�'޶�?x/l����Ϡ���n����w&�I/�_�l�1�y�A������kne�aR~^1X�E����|��_X㧃k=sM�_�����z�|��y �w�d�����cKv�����=]���9����eK�����,������M�}ͬ��@{���ϟ���r�w^�WL�x�&��Q?r+�%?d���T_�@�ӟ��/����q����2F���'����p��I�{�I����Z�|R�G�<���=�zd����������?	7_ҿ���_$�5��P��;R>�>��|�]��o>�]:��~���㏴ּ�`��>�пv^��Z���W����������g����9�9��ϳ�~���?+�?|��~��?E�oN���o��d���)�j� K�X�0��#�W����Ȫ�Ֆ.{��{�}~�}����qσ��nϓ�菢�j�[�^���l-?6~|OP�1��ܿ_R?�ǻP?��w}����|U��k�����>�����c����7$����){/�&?������
�s��/1������+�o�x�l���v���x�	`�J�í����!��>�o��6����ޡoO���55q�J����ߛ��'c�>l_��'��>���j���=��f]Y>_J�����%�Z�1���;��[�'Z���' >�ߡ�:��=\�r�X���G���XC����c�>5����z{i��_wE_���|������񔿆Ϥ���ߧ���FΫ��]�������:�kK�駌���4����1��L�s<d���Mܟ������쌿��b����������][Oe�kV���Z�#�5��5R~П������h����H����=����2�Y��<������yv�jɇi��[�C�EwcB?��zO�������k���A�n=ޑ����`�>߿�zEm}���ο���;�]���q��\��`��^^{w�,޶�c�����I�Q��6�3Q�K�����h�
��y_�i1�?�k͇�jm�I����_x�<�;����_�NA}�/����"���s�������b�}��x'�����W�y^���O������a���!�%��<<��qsib=����	����;a|NF�U��@ܶ����	>|߄�S���#����7�cY�U���%�k�/���L������O���^���g?������ڦ���Ob��<��xY����w#�,�Qc��M�s�&����_X�o�߷�GR^��⇔����n��x�@{�|��oy��o%<��&��e�]�u�~�������wy����O�_�/������Oc��Z緝>���l<���'�Oh�-D/�}�I���']|c��]��و���7�g�L��5���������Gq<ɟ��??k��}��@|)[�֡?Z;\���Ͼ^Q,�n����s���e	}����H����=5��}-�í�j�s�9�~�%�n��೑?�?�B��(߷ �����{�.ϵ����pQB/�#[�Izf��=���/�U���w��\v�K?�7L~%�~��?������Z���Gz�sM����W������5zd�,�k�w�z��3���#��_k��ވ�i�7������R�~��W�/{��sO���.+h?��j��?��f<"��o�s�8n��C��Z��{�{jw�.�T�ǣ(���;���9�A?���J��
�7�ͮO.l���/��/��Q����_����z�[��������߿ ��^����;�{"�/���`!���^�~q�v���??o�c8�^^��~З�L��������>��($��2����]�p�������?�Q].O4w�m���+h/o�j����z}�e|�;�a?���џ��қ�+��zY���AO���1��V��E����r���P�A{���E���b��x�.ӿ-������.1X��ϧi>��X���H�}'�7���w~P�}=����Oy���^�����,�P_g���r�F{���{!��{��W���+����L_H޹�و>�����}�?2��y��_�?��7�<�dk�����d߹�U������19>��Njm�4�/�Ə.��ǧ�}?� �����/�3�ߣ/�y��;�"��&3X�������=%��\�v��J���St�"�G�>���,��p_����_��-�3��ƛ�y=����C�k_%����z�>����@�����3���G���D�4���ɯ��O��=��yI�g:�O[�Ė��/�j��y���G_���q>�\E���+��,�$�D��k}���V�O���>�<_��~�4�6���e|�����Ɖ7�{����'\�'������H�E�>��.��+�/��-���~���5�ؾ���s�wVR��ߗ�ڗ�sy=���_���e�{���ۻ������F{\d��i��|>d�h�j0���(U�}
;���RH�������=�����@��?,Yr�����e�Ͽ�F=�q~��=��>�j����_����s��<����ͷ���	zIB?���"��:����[T�c�������f?�y�;V�������#t�N}��?����"�H�3>#[��!���_k	?�~*�W�G^�������|�/5��׿#����O��d����_>�g�/��j�׷k�����E�L��w��kng��l~����'����s6�~��{ў�S�GX?�!>�/��������s�f<��y��)�w��N{\�����x�^?��7b8?gp�V���A���W:�m8�=>��_�֫lO���N���?�O��g4������޾lU������������Fm|]>1��_���/�����kq[LȘ�z|�~�~ޛ���	,Y����u{�������y�>}������?7�^�?8�������՚���#I�ٗY���?��|w�(�~����b|�j����5{��+��g��k�N�O��x��ї5��姑�7�Oj���<�ך/�bh�<����j�������3>���_�!�ǫfOy��_<�@���Q�������Ȗ���k������y�3 ~�{9��+z���SО�1�t����oµ��x�A��@}���'�MK~n�_�Oo1��\/mO�k.�x��iѓ�O����?���w���S�OyG���h���o�����Ϗ���Y���`���G��2~a<	�����9�я/�͉�~���W#����?��<?���|{fR�/�y�=2}(y�m�/�W�?��vx�˅]��{�E�w�>��������b����U_�^\ҳ�L��%!}��}{v~�f>r���a���'?�K�h68?j���?�������.r��E��o��[Ύ8�-]���ȟ�o�Zoƣ	_���{�H�>��q2�뻿,}p}/\�_Lz�>3���oK?�iߵ�ǚ��1��}��ԫo�Q������>Z�3�����f�ףO���~#��~M_:}�^&oZ�tg�E�?��`�j�RR��r]�����lU����)�?��I�~���O��l�����}˛�o]��_�-��d�H|Z鳶���Wm�orY��������^VH��c����Z�wz�����n?�g�Fۋ
=yߑ��?OZ�w�}v���'�P�F�S<ח�{�5�����=�&�h����O{�.�>r}�#���������i�[P�L������)/��Z���D���u��i_���|g~�G��׷��s{}F+o�a���Hm~�_y���ᝠ��E�G���:��ץ~���=]��x����x֦���W�mr9�[��:�g�������$�����-{Nk�j�^~{���o~����G9�����+�W$������W����������ʻ=rr��3���Z�>�w|�_������s$��4�|�������Y�~_x6�O ~�?Wԡ�'�?_�/��=	}"����a�u�����_��n��t�7���唧6[uw�P�����?�����0�6�?��?�O%�����M������?�ϵ�����������p���_x���}��><��髰z��,���١��j�>�5ߓ�O��'Ƈ��S�>%�NG��W��&�?U��,����U��v�����E׷>�%O�=�o����f�ww�_�G])��-}o�Wv��
x����#܏\/Y�w���^{Y��x�l~)��7���$?���F����G���oC����^�#���/��_�g��A���V��4����_Y�{?�i��އ��,���!%O.F~ޟ������7�|�e^}Z�g���w�Q���L�#e����?c����_����+�����$�Z�_����e��L�_�j����c_���ߚ�<�·�_�I�,O}A������Kkя7�^e��j��ۯ����?�om�y>�����
��=������nzz��m1X����#��;��Vcx����~��H������;�Oc���Ί��!�H�畏�d��~�/ͣ�W��꺼�/�ף����Z���5���=�৕*\�K�]����֯�~�Yi�?R�7yO������Y��V��ez�Y������i��[.F_����=Ay�7����=��s?����������OF����(���C��/Y���R߳<ҧ�v}�-�^�N�7����}�7���o���?��:��I�����4?�>
��I}���/�b��e�_�\��6��i�w����!=ÿ�����Ǔ�n-�����	�_�?����?��O_F|/,���~+��d?��&�G���e1��:��G����?|�K}����	߃/G�<~;r{F{���|D���W��5������W�}=H������P����������O�v�@�� ?�^��������{c����i�W��l?��s`ꇵ��ײ���﯋��<�l+�/�����Eׯ�K�7�F�������#緾~���5����n/��fpM�9��Xݧ-����]�r��.Y�Z����b���`������·�����g�����E~_��#{�C�q����<���O�d��'���9�M {�	�!_�<����{��?3�IV_&?8_�Q�������ܿ(���iWd��#���3�/�6$K\���l<�"��O[�Cˇ�	|�#��������Ӄ�/WF�?!�=j���'�W��h��ϼ/�~�
��w�L�����o�ܞ����r}����7��/\|?[��[��W@?�/b8�����ز�_\U>Y�7B�y��%�����h��G�E��2�S�K����y^"[�R�o���3���M�#��=�{���?�����F�`һ5ҟOE��E#��ҳ9���Y�~���S�_s7����J{3�E��j�������&��FO��߭���)���������z�w|�jO��?�w�s����ί��r����U����m�_okm��ȶ������k���i?�<�� ���~���)�o���9?�������&����y�M&���#�Ƥ|M^x{5�R�~i������9��Q�������z|�WY?�j�]�ӫu�Hk=ݚ-�Y���5w��C����J��?�~����f�W��χW�S���3{^yM>N
�{��ūї��7�?3~3P������j���O ��_�����ʞ}Q��������׀���MEv�����O���ϡ�ǐ��p�_�t�0߳Z��~���g��������N��ّ�W���?��{"Ig<eM�d򒰾�~�����\����}4��/����|K?�b�����xJ1������/�oHO�����W���y���)k����s��hm=��O�=v��'���a���R]�לO�x䖿`y�������`�W�/�O���sҟ��^t|������~u{C���� ����O��g����󯫍�9�����>�5�=~��Jv�_{$/�/�|X��m�������]���?e��6;�����ў���>|(����qy�%�Mh�5]^�U���Z�^�������L����'�^�����+�D/ޝ�?���l���������*��}��{}5~����䟌?�_����{K6��񼦍����$��9~���#�c�#�����F�%�N~�y'��ѓ��'����@��O�~�[�I���W�'E|���慨�zQ����i_1?�Z�nF�m1�o��W�ߟ/���}k����s���m��*k������ߏA��}��}�]���B{Ao�П�3��S����6ė�mG���H��'/����߬�kv?�l��`���w��X?�#��b����a�_�ث��A_���k���x?Df?�Cyފ'��]1_��l�g��J�s�]���1ܯr��V��0�ϗ�������.�w�P~��t�S����<~���O\H�ޗ�%���;ȟ�!���do_1���K�4��L�k~�� ^]C{<o����q��3�A�?��/^{���`�`�'Pk/�?5�ڲZ�{�����2�g������������N���ϼ���'��W�/�)O���<�E|4W<�wG�	�_�O���3S����?+[�-s��Ӆ�s����<�K��� ~��&ɿ�%���i���\�2]�=��в�~.��[����]]~�q�Qy{{bO��_
tg�x��z�x���Ϸ<+)/{�폖>�����"��{_-���׻��8����|��J{N������n�j�����%/���-���h��&��q����Bm<���F��=}=��]ine�./�����$������\+�IkG�o��-~��em~{{����ߗȃ�`I����4xO���m�O��]�-�̟��U�EK�O��q<����}ꞟ�Q�>��Io��{߅���Ϥ�k<��"}���GX���o/b_�ٿ��KfoʞXK�A����F{�Oy}}#Y��I�������1p��m��Y�>?��t/��7.]���끨��p�9�k�k�����(�W����)�������ў�/�7b���z��M����^���$����oA��L}w�����w�k�/��3޻�_ޅ���;�?��d�WQ����R�I���蟒�y��>Η�6���
��!���n?�on?��]�ߖ�?�������W�/��P,��W��}�Y;����>���䷿����'��/��ԗ�^^c��Fu���/���u�M��s�~9���_��ެ�W:A~_ҷe߈�Fy�_��x2��Q�w���OZ����s�W��sk��Y?�|x���})��G��/|i��c�?���'�O�\�΃���O�E�~ۋ��ߌ>�6��~�n��}{dw�������'#}���G}1��/�'n�'�F�gE~�m.�ϵR�����Z/C����� �K�ח�g�w��Iy����R?����ʊ�*=_M|��Hoڃ�诿8���|OX���$_���1�/�����ch��qz���[?/�N�}���Mko����>���<���뻨������l��n��M����c����5���?�����ьG3}�����|�}n��>jɎ3P������ߥ[ܞZ��}�o�D�:V~�����x"��%�/w���T8����񀔯^�ʾ姍��+�s�P�����ƫ8��>������J��E�}u��No��8���.�
�9>�/%�����v|YDN_���Z;O��|�'&�"�-��O�������[/?�<��=�.����0�o��Ή��l�3�O�x���W_��Z�<�4�	�����ޛF_����c��i���%��YK�g{���l�:��E$.2����_r|.����?d����}{��E�t� ��o!����>^3Y<�����_<\~߉�:����+��A:�5�y�_�����Z�{*���k-�(�O����e�p�������O�g�Y��+~h�￫�����/z�=�L���Qy]�?��ׯ�0���s
�}��{zҞ�=^Wk�ϗ��6~�j��Eҿu_㑅�Ǔ�����������sk=#�OAϣ��;�o쀯x��$k�������o/��}��W����k��~�1y���KɊ���ć�A��=�����gu�x�}������I1��d�d�{�����E�G~by�w���x�-���}}���9��1���~p�|�~�4�/�u�?j����G�\������:����$��o�WR_˾`~���W�SP����'��L���^~��?��C{>���_?�#{���߭��l������.�k�?//|�"~����v1����㤷����s���~�?��}�0^���������m���F��+��*��5>�Q_�P���|v^����Qڇ-{S��f�d��S>s^s�O��D�u��?�������x�w�B�=y>����Oy��D��F���o�!?e�k�����m	�����>���r�_���v|��O{]������$~y!�w~�C��z��a���#�w�!������$��Z�\/펜�Ho�7�c�?��_/��Kz�6�gzC{��g�\?
v��y|Ǘ�q�x_B����yL�'���I��Om������q����:߲-��nɻ�{��%�/-��J�3��7�g6[�M?1+���_����%OX�ҩ_<?�O�|F��7���^�{k����,�Eo�?����|�x����NF:��S����$y_��w(���������@<E����so����wƐ2�/�(���������4�����I����d�>�zy%���t��My�x�����Z8�ԯ�_���>�Kb||��0�r�k��I�2�s���}��gm�9���vԗ��V�ߊ�`�~Đ�ox��׿O�~?E{��� ���j����z���i�w���=����������e��ޯ�[v�Ws���g�!^��{�x��3�/���p��v^���_��a>�қpm�+��I����\y@��o�~�Ӳ�����EzQ�О����g6��_��Zt_����~��YK�%�Z��dP�?�g3����Sm?��Ӹ>�=��,w#�H֗ɯY[3��_�b�D���y�V{�.E�~Y��#��5V~���CT��Q��Ӽ?G����������}bx>����#�����n9n��������x��o�h�[�+�3C�8�_���]�/Z��N��b�>��m����|{��kWZv>��	p����j���oޗ1N��1?�g����f���?�����`�g���� Y�Q�5?|���c	~j?�?C~n����ó��6����xg�'�X�Cyҟ��y�9��G���Gg�kny�e߬���WD~��~wK�-{H���J2�V���'G�R]�~��d&c���婿N�|���>ǫ%�j�Iz�}����?l�����_��|���L�Wy����'e�/��r���H��n�~�_p�tқ�탐��W��n���?e�y��x��w|t~�����S5ޟO���G��G��˷��y:bh�{~ɖ��/�+ȿ���>m���W��W�Wd��'X:ϓq��U?�)�=h�c������$�<�H���$�5�O~���7�Ϛ>w����Wj��3���T���tV���p}P���]���`�O�_\�j���98�䏍�+����򚛙?P�_�h�����@Oޯ;#�)O|}-�����O�{���%�菟�w���w�9b���
�ӟ��:\��r��c:��j��>������o�}��_��ztRl�M.�E�/'~ҧY�	޷�O�������Oy�%滟�����ck�h{���M1ܯ�~!�������>ښ���N�>������^���q�7�|�ޙ֣~~Ns��d�H5������|�����7��m�������q���w�����Ҳ�J���%���	��,U�����d�5�d?~ �9d����џ ��A �����/ǫ6���*o_�ˌ�s�K����W�?j�Ӂ���R��׺O��	��NѶϽ>�u�@�^���7���UП����������iݯ��������'���Gz��S�̿-�����_h�O}q8��r�Y|����(�%��lp�o_u�֓��\�f�{f����c���_�g��_/3X�[K���Y ?�:~����?l����l�z�Β<�W �|�����h��p����%��=}�I�5I���Y|�x!;O�?_���_������x���A���ӷGߟG�Fk	?�(Z��!{����K���g�̿��PP�'�w{m�	�Ώ�����E�c!������ |$iO���;�[�S��}�̟�3���P>s�g�Q�#?;?J�5������?����ހ�l?�&o��E�u��^�l�k樏�T����3��/X���0���C�����e��&�<��^ї�]����;��g��ʺ�~!��������ш�������z<�V}|ϼV��&o?*�����������5~�����̿�4��d&�]^���+���Z����]�~��=�Z�I}��L_D��O3�����i_�����C������������n���(?�ח�[$kn �<���g�}|?��WYƗoC�+K^����0���ߕ�?9?hl���P6�?�p���M|��>��nw��h���[b(�2���ɀ��ҟ�_������^��Ax��u�.�#������,Y�'+����/-%�i�G�w�;�K_>8�_GP�?�g��Xǭ�t����E�ݺO��������K�����s�By��Gy�(�=�����O���j�����i,}��)���p�����w3�[���/����W~����0�r���S�o��C�H~�����շ�ǅ%_��,��pm~z��kQ��Z�������m�1���t��h}�`���el{�A�{���������'�7�����_���V�����j����_����q�t��W���w��)����S��^��~�E��>��,������>��P�����ד�m|?���'ύqzp=4�ec���^���_'ޤ�OxW��'�j���kI�����q�9=�{�u��|�b|��_>_H�#��/\����Mw�ײ9����1~��~���_XY�.xz��s~�x���Q���N�m�~�����e+���������g�-�Q��~�,Yk)�'5���;߇���=b���}�=}#R�;�����q���'b�ol�a}%�����>����~�_-?��g���ٿ�����߇����=�u�VlЯ���?j��}p�m:�'Ͻ�Y����&�f3�D�O,~~r�_�#�o/����!��奛/���x}�C�ݞc��OE�uoC��s�����΍�>�}}\l��	�{}���߈�|����ߚ��`����?�O�������G��__J�>��[K�M���|��~�/o��*�/E_��w���K���E?_#�*�O՟��/)�?����o���~yf��oUY�?��#l��}v��~^P���'׻�WPv}s���Ǒ��?��U�><�Qz+���1���x��|��������]��'�>O��g���<��W��5����'}���(��k�l��m�G�^��lv��F�������G��M��O�_���|Ri�_����7��}v�Q�����f��>/(����#���?���<S����W>�������bf����Y�����/�!�Ws��Se�K�?}_�����M���G|��N�_����_���E���}�%��� ꣣��_-z���O�G�~�?e����F�}A��_�[���"���pw�r$���p�ҟ��Џ�Y��ѿ?�e�Ivq}�Ż���V߶b{���-��[Mb(O������ܻע�;�=����^�ʺ���E|i?�����m>�1~���A�>p��xz�N�~��)��WD��Ǉ�%��?�G�=G��|�E|X^k_�߳��<���ߓ��Z�������ko��7��Q����O�]=OE�._�? �55X���s���_�E�������W��?��׹�.�}g��Ǳ�,Z�zi#���d��<�����?�W�7EH��<OO���k%���,G�?�ז��d�c_%�����}C�����l�g�o)���Ö��|]R��_��k	}g����O��Y���������0�c����E��u�	�/^��ď���-�}��;@�3�W~߯��-}�x�3��d?`��*��*���,~��_�j���?�������=��k�/����>�x����G��XR_Đ_����;=�o|<���z��1�~뾎��*�c��qH��	�'�Uu��`�+�y���G������h�J������>.�iB���s���M�?^<������$��>r�d;��xQ��[���0ۿk�[.�����Ô������P���҃Kv?_E|hO1~�竹���[���_����%���?����9h����+���㡿,�^c���2�[�|���p��k�s�
�ݾ���o1�^ _�ҧ����;��`����F�����|���M������o�F����Y�=�b<x� �7����AM?����e/}&��S?�o��8�����}8~��q����_q~�DW����#�t��:�[�\��xy~��o@��}_���1�g��Sy����@��{���"��m�oM{������&���3|���?�����B}*���W����Fy�7��>H_�ė���3�s)�X~_�N�a���-��ew�~�-��F�������Y	="���;���п7B���x��bl~��ϊ��i���<ߓ�^��F��rԗ�Q���K+����5:;�����޻�,�9�?���K�/ǫ�_�����˥�����Cy�7���|Z��E�s�y}-}��\��@{|?�����}M^g�������|<dO݂�����5�����x?�Mv^����~��	�\�k�.A:�{��v^t�R�r}���|qy���q��/�󬍱��<�-�/����~��:\�oN?�N�?;+��my���@{��,E.Fz��m���e�~��e��]8�R����-]������R���q�����k���q�Q^0^��䧚=E~��>^��M�c�;O�����q�����Q������yI�����/�q�/;�zF��^�|�������k��������햲�>�:����яG}|�0~/���>��>�����+v,��<����_����_,�#Hw�Uyy>2���"=į?����$���������&�+&1^���/K���΢O{�l����
��`͵��-�'ڵ�����@t>�7稯?��	��b�x}ڷ��_oO�ϋV�l��{o��~��ϟ+c|<��ߌf�O��{}�c����~�R?d0ϳ��qX�1\�s?��=��&f}�����>��\V>����v-�/b�� ��%1>^l��iOJ��<�>��J�eG@��a8�j���	����'~��}��/�������?d��޴���l�L����0���X~?��Z��=�U������Iz��W�&�����K�� �3�P+���菏������U��~�)�-�9H�#��e�f|�t�{>���⯏q���I�my~���Γ�=(�{��3�C�,�w��[v6����9��}F�?���d�������/�>���.������Qƿ��,�_����g�C{3 g񺬏�����'�O��m�G�/�G�߼��pR~��J��㣻�n���e��t�c���➿����$}�.��h��Q��f�����ڊ����Y�9N������/>�����?��N��ѷ_�����5�N��|r�d����a�D ������g���e���F��7������;)r��?xiv�����1��-���I��;`0�V���Z��d����#c|��$~��{kI}���B����/⍗��~�s} �0~�C}o0��%���������I�ӟ���ƃ��h�d���Ϡ~��kM0������g�흇�����?��x}6��4rp�>����+�{R��\�|���яTl��K��������J��/���sk=��K��yާ����oк�����}e����o?X��������x����x8)^���D�d>tU���/�W��e�_Z/�yʃ)�S��~��?"�?y�I�_��������{[����C�/S�O~��/�<��7�;ϳ�t0��vE�~X�OɆ�>�����쿕Џ��.��l�D���U]�zJ���ʃǗ*�_1���"=;��/�m�G��E�>B�X1����"�����<?����� ҝ��Z�O����u��+����ď�q|h�Tqy#�<�=�L'�ߐ�{��������~���?��#�c����E5�l�+=�����l����.��l_���/�k�38~�������>*���/¼o��ǻbh?x���k�&���|>K9���W���O�7��w���y?2�����=�O������y�������)����xB�G����;c����!��_I{�������7�i��[[�1���O|&	,���H/�!��~ށ�4����<����|���u_��M�������.ώ�ϲ��k��4�[I�����9NGy�/��$��W�&��}�Wk~NP������3n�����������!�����S�?��U�7�y�Q���4>�-u-�񻼀���K����x���O�����?�[�q{��c�����ޥ}@|�^��e��W��a��(��#�W˟���sY�N�&O��=g8g�1[O�̯?��~���#~Jߓ�����dzF/���1.�p��l>h��g|�����6X�CI}���J�N������wX���"=�ol���Z�?xy�����P���ڏ����4���e���c|�����U�d�����ޖ�_C��'����?I�_�'[��$��y���4����?�����@������Hz�7o0�̒��[��o>cp���C��bקY<z��2y~$��g�>/���y2����+Ϝ�v^����/ld}��Ӛ~�z����/d���nM�S����������������/�h���Y<D�~_K�\���=v��a�3�i�/��qD���=����w��}���������#�?�?���v��E��O��>�[���x6�W]�����迏��p�_Z�������8��p�����y�Z���߉�����s^��D_߯��]��Y���� �����L��i��Z&Ho�/��8������s{[}e����d�߷*ۅ���/��?����A�����c���/���a����i���^���I���YC��|n���b�8˳}��ނ�k��>��+ȯ�Z�W�ߟ�l�<s�)��п�����/�����]m�a����菗���_�П���C{����y1�o�}�S������bv�C�����c���?��_"�oo��鹯R־h���������$������<�OY_d��*��R�Ӡgv_�b�����/���ƛ�}��y�=��?q=�������o�K"���M������}y?<�ӽ�B���vw������Ǚ	�����'�t�����7�|��~&�?�j�?�e?�q�?�zKs���!��7�,)_[�y{�ZH��1N_髧L��Zs�i|���"�/2z��=ʏ,�l_?oN~��[��yE�7��y/�g�}��<]�^��/�>�O���a�^�f0��I�� ���g���5�j�ALP��O����|�|�������|$�Ǘ�騮� ���p�����#��9�/��of��W��i�?�=����D���/�O�oL����}[���'������[�gO���¯�U��&������)��П���?�b�������e��k��|�y���*���W}��k72_��#���4��;��������l?��;� K���P���i�S�`�����J��U}=��C�g��-��+���&WE��k�s���;������}�/[:�E?��e�Wc��$�fO9�������xg�zA����WJu��Ym|�ߏ���������y��t����A��ӧ+�ٖ�����}�޾��{�?K��~�l��3X���w|�[���G�H�zQ��'�#�?ozV��a���Y�o~\Ob�5~��3[�~ �}�l��)ηI���������>~7iOu?-I���:Z~/7Xs�Z��[���������b���o�`�_�z��ݻ�e������|�}W�s�StW�d�o��xލ���W��>���C�e���W�3�o9�OXk�o3���{7�Պw��j��S��|��R�5�%Oy>��k���
7�o�ޅ��$�����'g�]���z�eO�?Z��{b��\�M������bߥ�����V�|OR>b��C���'��=������ѷgy��������o��x��������zd�Z��ݏ�~�����G�<:㳻�_}Y��Ozk�}=��4���+�K�W������G��+��{����oH�G��O��{\��=��p~X~�t�=�A����^��1ԧ=e�z���.����������4�����g���x�|����Z}ې��a��w���g�il���r�������4��b������B��Z���A�>k��x���/3X�"�GŦz�����G�g�8���cXO���.�$?�e�� ���(�ur�`�He�A�,~��������֧�
I�gR�ZܶFv~��g�Y#rCk��{_Z>W���{��=�o+��������t���B{O�C}��[��$�ԇZK\o0�O3��ߢ�þ3��?�z���y�����Ê��}.���nO�>C��џ��x&���w���ߛ���r���_����ٟ=�_��Y�׹|�`��F��F�?$�>�t�����������ΔG��f}�+�޺ϐ�Zz��R��QY-�<�o��(O{�gc||[�ɏ���)��1}}��-Ի��u1������ߎ����Om}N8[_K_�%��Y<bT���f�C���F�l�B|��']����y�J����A��mȿ��3����������u��!�_X�|�����|D<'���_m?c�x�i��(ʻ���k������D�_2�����?�uE��z�뵕��{���>���;{?k�__����$�KzR�?�/��1�<�|b|%�M�|k�'�������t��>G�	K7�x����~����gc6�~�}�>����_n-��џb�M>�����?���w����r~%��F����ߗ#ڸ|;=��\����6Y���7t���pWd�&�_o폷�i ����K��ߟ"=���[��ȏ|�@������*���~{P��ЫȖ����8��W_����>�I�l�f�:���O�#���4�[���i̷<�\���~���_(_��K~����?+�uy!Z�y�{G�|�~��"p���Ƴe�Oh�p}+�s�Q��>�{����q{Hs����M_�>�?�����I�Y������o�?&\ӿ���t�3Q>��\��E��� �����5���L�����c:��;۟DN?���E�����Ŵ�͟�1�/��`�-�_����F��T��>��"�����w�`�3f2��9�)/��;�w���$�О���<��SW��k������Ǻ���lK�W��?���;��@ٚ��䯝G��m/D|"��#�7�1\y����&���ByZ/O߉t�CyW�Z�xa�;���N�}������k�h5��<�*���Wɒ'�8>���$��CXk�G��d�i���b/~�`�����l_���f���
���O�A���}D<O5�q3�ѥ���~��&��'#����Ծ�З��z}��=��t��9��G�����睺�����I������뻊��o���1>����_�����~.�]�?�}�������[߲v��{T�W�>�����s*�gy�������C4�.�4vנ�I�K�EO�W�?([�_�5;�޲ϙ7�w�ϻ��e.t~�r�CNO�/�L�"�}�c�(�O֟�\�)֊�	�S�>�{&��^���ݟu�T�Aԗ�/n�����������:��Y[c�?#�����E�כ�>�n��z������<�|ס}��F��w[��+R^������"�'�1���?�#"�����}��+�e?NѾ�+z�}�D���Q]�	�e�d�QD~^�bOuW"���������7IW��铥�F~��U1>~�
�q�ŋ.�o�Q��I���7����Ϗ"�_��MhO�6W'�_�xɖ�x��6�2��y	__O��<��_>��/���Do�_k�>m��O��7�-�_�~��)����~ޏ��S��D~������i�P�G�����Q�l���ׯ�3�^�����(_��5=���i��ܾ؏��ye�]>��\����g�ȼ�/�K��}J|&��g�^qX}�}�᫯�wg2ad>O^^X�/@��������[0�-���$}^X�q����G�O����e�f�/��%�����@��/���N��������ڿ�~��7���B_��������������g4������������z�g��������'�_�`�Yyֿ��M�M>>:K��ﯾ� ��p��ߺO������e�{���SM��|}i���'k��IR_�%���j�{���O2��h�c�x?�|�x
���Pߜ���|�5Io�����.�|<���F�;?��~���G����h�����o�'��{sR?�Sޏ��������皟�~��9�G����{��ͯ������#��?ߒ�ܿ��x�П������^@~����W���sZ��e�I��]��i�oD�Oҕ�7X�u��<�M�e,�㗽�P�,���<�<X5����������Z��u:G�M�/ǣv�c�S������N|�]��W����S�>l���� �Z�b^���?���X�y?�O-�y9�7S�?����_����_����҄�+�.����?h_��:�OO���c���P>�?���^�����zE�>�����ҩ�{������G����>+����Y<��:�/g����9}Z��<�Ъ��E�/c���y��O��I��%�����|v���B~�y~�˻#������5��_>^�Ѿ߹�O�>:�'���&ԟ�7���姀�c��oğ��؇#/��~p�����樿��};�?B?��no1~Iy�x������q���'о��=/_�G$����U��?(���szkl���[��{>����Y�3߇f�Ӄ�Q�'�{�>ϣe�H��^����<�!��g��tz�{6��`���{����V�w{�4��)�/�;�Gc���_+��'�����U�N�f/;Ҟo�j�����6�GIk�J���(���y���d;�����k<�3X��ϋ��|���_/$����}K��#�����O/U��|&�g�t�˒���}C�w�� ���(�r����|n��%�� ����27�SY�����}��b�h}$����⿫��y@�-~����}�:�����F�`�2a��9�������s�S�O��RߑV�ֆ���ɝ��%�����9r�N�$�/���g<����/�=���'>_��>�o{�o$p��{��K1�?W�e��P�2}Cy��6O1X{�~���/W�ߗQ�\������E?�J���Ї��������_�O�߫�,�k�w�E�>�]���4�.?�Y��E}<���3ަ�>ϓ3^�#�ono�|�_����|-/6X}�x�gk�W$۟�������7&������Iµ���W��>����L?i���,��3�ߚ�ꛯ'[�J�<��{2��(��Y�ם���^�������tyf�����x]\�w)�O}}*���l_{I�0X�����c��֒����w�p}���~����D�����X>��<��.�ӟ^;�I��z�ǃ��ظ��x�����>�������z��C����k�2.�멯h_џ��Z�7��Dz?��r��o���%��Z���/ݖ�&�m=5ym?/��c��<���o��A����������� ��.O对!�ϴ��������}��ۅ������|e�?�?ׯ��,~|8�{������5�5xK�7^߾��x�)����<�G�����k��?��U�/S� ��w6�f}�?���k�q<�?_��Is>����}?��y&Í���y���o�ԯ�Q�� �Q|>�����3yN��L�������m��]��ό������g�ҿ	�g�@ګ��=��y��z_}B�.�~�џ��F�;-�拏<�R��¥����Gy����?�=M���շ̿���K���\��?��7Z����M�_��W�1�s���Q�1x�a���7�??ɿ��Ok|(oj���;���{�xޭ̥���ѿ�2g���O�����0����F_~�޸��<ϳ;>ڟ����w�?K���Om}�����Gy0���3�W|8�����g������p'Y�	�'���(���G����yK/���oB�|���C���w��SK��ֳ���@}ˀ)?]�3������oE�ܚ�_~��{>�c|Df?H��JB_�']�Z��k�Iy���AO߅��E�?k�]9=T��}i�f�Cg�ĜO�������Hw|4��h/b�Y��j�#�������y6���3bx_��'}q(�㛵O�#Y{���W��? �="��z ?���!Է�������֒���>��$?�����[9�O#���y�9k�K�o��/������~�|�e�h��֢;�/���'�K���ֶ�_܃�<���������{�\�q���4��V�wD~oٚ��S_�7v{�ӥ�5/!�b�?b����7�OSk�N�_��f| σ�/i_����Z��ߌ�>���t����z%�/`�]��{�onO��~�Im�z��!~\�ii��'%��J��������k-��P��G��x���Ǿ$����o�ޏ@���+��~ߓx��C���ݞT]�{��G�;%���ZO��s=��b��ע'��@{��ߒԧ�e�g���1���>���Y�o�>�;x�1�c��	��;|=}U���5����_J{�Q���9?�~j��,���j����r鯼�^�l�~�gy��A~������󾜏�#�_O"��&?3�ſ��G��yj���~�}_�?�y�F���?��7�y��w�3���%t{q1���%+x>�ۗ~��~�?��f�q�#�u}��%�:���8���I����>������v��m������ӓ�������9>�[>ߟ䗽�x�7�ג�������������w�M:��_oOy��Rp�������n���x7�G�+�?>��2�xIV�=� ���zS�jo��H_���9�k~Es3�_�=���O\��D?�P���#=)�E�5���ya}}�-[�f�5�_]��|�|d�W ����%�k�Y��EV��]y��͈�z�������
�OP���+�_k�O,}��j�G\����ύ����{y�˔O5y�o�`�ߜ󭷟_�S�>��LR�㯔���~q|5���q�%o�!�_����}�O$�)�)�P_wKA�W�����G~�Y���i��x����Cm{|.������'�_��U��\����n�J�y<3�I�q����s�G�yɪ'��Y|�R�� �4�������z�e��~V���?���з�>�=�������~wk��h����#�k��3z��'K��c��=�m_���_y?�ǭ��/����h��Rd�����<$|r�]�� ~��,oE����Z����'���nF}>߅�ۛ��~�H��=.x������1���d����n����6��{na�/%��~`����${�~�V����I���n��}�'׷��Ry���g�����h�������gY�t����|}�_������}��E�>�S���p}��%��|S�}�`���|k�{�Ox6�N�g4���g��V���v��+S��Cc��y�Ǚ���_.m������[�����g+1��r���^8!��ٜ������|�Ni��w|D����_���s?�~˱q���E)oy>��VV?ﳉ����W?[�}���]����Y���ێ�Z�����^+(��-��o��~�,����4���'�v~9}}GzI~���=*^=����xA�{��^��k��h?P����G��\�Џ0����랜������_ъ�%��c��'x_���Z���,5��?��˖=5��Ͽ�I�d�>/�O}]G�����O���x�E�g|*�z�q���ɷ5�����Ϭ�������Z{�O������Y���g˞d}�珍���Z���??�Y����>�>����������Tl�?\���3ާ%�r�ryC�����㥷P�O�%\������]�'�O��������_�9�t����Om��S�p-���>��xߣ��~�h��Oj���5~�L�O����1�w�����Gk��Cy4A}W#��F>���ǏoD^��O_?h�^���񧼑.���5>.4�OJ��xt�D?>��}��>e�E��"�+~�|q�q2�k�����o�Z�5�ί��<_��������������x%Ͽ�?'ly?�l৹��Tw��y�3A�i����q�E��W_���ߩ?8?���R�uI}7��������(�������<^��u{��7�/��-�ow�U�C����F�Y~��}�5���ވ?)�w�> ~�Oc��_�P^f�'���`��V���6?��]���H�c�/���SP^iǒ����,M��{i��2�����Ok����>�����%�>c||��=���?�|�F<Ey����F��u�����$�i�	�ė�3]���+��������bx���&�ߤ}�گ��W��"}��7^���`|$���d�}�?���J��+���#}j�Q��߫�=���j���5��������(����ڢ�i1�ם������?!���ū��-|���o���}S��l���{}���U��Ow}�\)�����lB���j��K?P��<�%K�����)O%�}W����Py��?��֨��)�s��c<�-���k����P���QP�*����;d?�`�֪��On?ѾR���D�>�_�'!����_�W%�i�Z[��q������h�5��n��~��?��y|DM^�>�̾��U��K���%���-���Cy_���<����?d���?���U�w���Qi./��KP���i������~�^T��~��/0X����ο�W�s~�}��?�G[�9���}�O�۫��L��d�ɇ����+������������D.5W�L�����|���ҲxWц��<���K6�������������<T�|��+�ov��Q�ǯ�~��x���W���x�U����s����w�(U.������a<���I��P_����̿������t�N/�����>���K:?��q�6���W������/z�����ݫ�������qy\�0���#���-2^����'�/$�z��@Nψ�x��_$難/�u_'���t�2��}��=vR�S��oO�|�������7��G��=���x������ſ��|c!�'���٨���ߚ�8}���U�5�*���߮_�M�)s��>`��&����H��Q��7�_���+}�|���X�����3���ʖ����>�?���͑�'�9��Ʌޝ�wz\A���z�=��������o�x�=���==���g�v�x0Η�1�/��#�e�6�>s~��ʻ���ҟ�@{*���w��򺽢�i��	^�}e�/��t��[����*�s~�\��I8����V{� �܏��xԥo�v�J��_+�I�����6����z�R���;}����s��1�"[�s���C{��OF���&_��pK4詹��d�����7��/�������Ns��<�����b����F_^��t���;C��wS������?ݟ�߂9�T��'G�����b����#�}UL����]���#��Ò�7!�����)�]��G?�H�O�9_f�v�k�g���5��? g���zk�]i/���/}��GN#�g�������c;�O�����\�. }���`�ov�ݜ��O�����������O�D��?T����i,/A{_��|�5?�~;}}��v�R˟U��d�L��=k~��^�����<���}o�߻m�o�S>��`<�Y�/;����d`&�V��_Z��qzH���;̿͝��%[�F�2�=y~A���C
�}��|b�bx���k���\v~@����/۔��;��h�������7��_���J��/ǌ��vږ���֎W��5��4��������9���:�AX�}��t���pF��#����"�>��?����e���W�?�֋>��J�O%��Vz�~�����t}P[��>�l%�����;!��?A���:�e;=$.D�Lҵ_�C��-��|��,�d�ww"?���#�������-ދo`���.?o��A�>ԗ�I�	��Ϧ����]��z��	/F_�ʷ����/6�]Y�wY|+�������+Y15����!1޾���/�}K<ހ��_�ğ���0����`~�u=���xӾ��=�D~�K���WܟE��h�6����޾^x�����*�x��HO�/^q�$�j�9Ο��������c���#�����/�~���Ek�G)���k���!���\�)�1N��}S�z��އ����8�L?-��.��x�i�O��sM~��ݟ��8����h��5���-���ʺ�+�ߺ��E��i=��Y{��|��I����m�_%���)k㳔�KyG|�v���9���6��yN���c�GP�5q�Q_�Wc��2����l����@ҧ&��0����k�[l_>��noj,��c	=���$?���὇ק�����a�> �Y|���(���X�G�}��z\��7�?����y>��m���x?��2~��/�~-���\�0�Fs��7�����!~�-����A���I��<�~�tޯЪ���YEo�Y�M(�����A/��lG�g��r�O��K�� �|���l�I���|���7��)�sZ���肉�)��?��n�_a]����t����W�>�#f�a��7���	��	�O�M�o���鬨�?�����L)�G��������v1<�����C,��\���$y�Z�/�釓�j��C��p��_���O�������ї��_�_�k�t��˺2^~������,{��3i�~�<���wYh�{�������4��5�D�_d��}��=�O�Aя����������`�"�_��Z,�8��S��};��o��;�'ߺ����g��l=Dz˗p��ܟ�_�;�1z��f�	��&��C˾tړA��K�~_AY�u���E��d��W�����KH�}�3����ѷG��yғ��틐N~��$n���e��,G�_�5m�7{o!P��S�?�wH�Y<�����![��g'�P�>���������/�����ZOR�~�W��O~֗��3���-����oc|��h�y�boM.C~�/����� �����#|<5֌�b[�D�t��?�C~�����}?���x�	�'��?�e�����e���l��/��Ț������w�Gݴt/�Wj�	���I?O�}��f��2��#)/��4��ڣ���C�J{��k�w��G����hn�<r��Ƌ��ы�� �Z�V|��Iy�g�����y�x��C���c�o�^i�x�e3^�����]�OAy�C8��>e�ϡ�ϻ��ُ�~����ʶE�_������/��ୠ��#���/��$�����</2��������w�����~��kѿ������w��ϥK>��S��{���"__�$[\ߊ���;Ƨ+���9�}�@���MΗ�<�<��)��|���o��g�0�'��^��-x�����j����/�}��Z���?���w��rWkA��T����/�����5���k���/%��|Y���D���F./[0��y�/�^M_s�C���a������D�,}��j����G{A�=�A���D��1�������)��o�o'�w�^�F?�ƒ���e��.�o���3���O�l�O���Gzo����N~�Z���zq."߯�/��z{�#��P>H���Eo�����KD�^�G�b|���l�,{(;���}~h��&�P~�x��˧���Y���>/��|��X���r>e��|Y�^�o��#�#j���/�"W�����I~�z
���ߺ���_HX�����_nOI���]�����1�D_���	=��w~�A�<������˳ԯ�(�W�ѧ�q�r?��g�滟�����f��/���Z�������ǉ��{v_����|=�_'z?:�������_ߏ���<��#&1N_��o�~�	���h_��]}��0ڛ�E?���(������x��?��+/2X���)w�a|��W(mj�d����o����F���0����
L�4�W�m?��T���������}��z�pM�d�/G�-z�G�o_�>�OmT����������a}�խ�_Z���E{[�M
�6?���2������/���jz���)x~���3��~!?ߣ�� ���x��y�g����{�l���k�U���G��1^��M����S���D��(���`�NӤ<��|�ѓ��������n]i}���u�:��^�����/�����_�w�_�~�_��/�ţ����<�⃘>��<���E����tV��m���d�߿F�M�^=�;0X���6X��������|�EO����l~��Fy%�w�1�������h��'���t��W�&ƃy}ҝ>?���������K���)?�á�����Z��%�F�P�?��?��0�H�ݑ��'xuj�t��w���{�>����������6������=��������~������^��^��=���I:��x����8�|��������hq�`�������YK���JB/���=����OB���iwW����|��}�+�GF�M��/'?��3�t�[�����	���ϙHg~�O�v�)�����2oΟ�?��)��������v|F��a|�F���+������𹨏��bx?=��N_�+�F��_�ou���%����%G���5>�����������'��~b<�b�h�e�ۥ��O}�=��u����x������|����c�?��+�,Z�?Si����'��Ɍ����gSL*�3�����������>�|���)�5����)�K��Lݷ��5�7�O��`�'����b��.��K�~�o���H�k._��?��������g<2�E���������|�?<O���ˏ��돈�����.��ɳ;#������?1X����N�����-���O���l���w�~�`��HO��?i~��x�
�`�/O�~�����/��.��,�%��|�,m?-��2[���M|T�ӏ�L�|S���o���O�`}]~J7�������B�.����Q0�����$�����J���cя�����,d������0��9�o|��sf��?zsi����~���sΏ�q|4v�?���ڭ�D/�_��Y3X���K�=ʻ����[���{��_ү5k��=]�����Q;���$�B}�O�x�~t���M�����!�׊�r���U����_��n���������"=;OFy��$���j�N�j�Q�/\?g���n�#^���(e;�O�/��O����������?�e=+IW�~��d�ۿ����7��y6�C%;n��x��@&�h�HV�zd���t����˟���1�gV^��|�&��+k�����<��u��t�2�_�}��+���ۓ�t�x��ρ�{%�����|[����<؟ԇ��-���W�>K�?K�$_��p���R�ܟ�x�ˢ�/W��|0��`����#�zk�.����y_4��ח��L��~�=,��V�[�[�}�d��`���yVf˶�2��[�wH{��q���O��O-�&�x��z����ҝ�Nʫ��X��<d�C���c�?+����鴇j�=�oY���j����ں��>Vl�Zҿ���k=�/}��Ĕ��s�z��{��?����i	��ӯO�^��͇N�����%���O��I~���oe~���ӧ|���z��/���O͵�I~�[��]>-?��|uy0�����^^F:�C�o)��U�:l��n��1�/���G����^��O,���~� �7�����&b�ğ�G�?~��b�1���/����?�/�����q�����{�!^�+���9�_1����*�
��0�����a?tg�[��%���z��Mǟ��`��d�Lv��p~�}��Q���P�o��/�8��_>.�e��Z����+I���L�<q�B�<��R�c��[���f��b��4A��sz��U>^\>�0x�qyB{�v>#��a�WG�>��3,��q���9?X~��-���0׫����]����I{������,{������&���,��K��P8=���������R�e�W2�i�3Xo!��H�p}Z��3������~�/ϫg�i����$/���QYou�����5����ov��k�5_�~���gG����q������>�K����T�|=/ܜ߸^&~��菗�ɮA~�Sҟ��GA��>��o����}���&h�z}�]>S���<��c�3}��=�C���L�����%ݟt��!���w��0>�˯�p����������Tu����5���s�:�B_�g%}{_g�:����eT�y�����/��1>�>L�;��߉������o-��A�⧑�������`�����|�/ ~�����[�I������O}	�g��^�+�����Z��OZ�d���5v�*��q1�~M���	�\>d�R��Z���P�:/�4����~Ei��WH6��P�Yv�����<���Az]��Ə���)�����>�������^~>D�o_���;[����� ��W���Aɷ��.��D�|��5���xo_��K/Fn/E�5�O����	��/�_�켫d���>��l�/f�/|o���a���W�o?��6"o3yԊ�}����5�a���W�ϥh��K,���~�Ӣ�O�/?Z�t~�>���d��?�'g%�k�!Z���?T>�F����W;/�����g~�7���#}�Г�h���t��V[����Vp��������������;�K!��<�K����CI}���pU��C����}E�d�K��ǿH��E��x�V�[���� �2`��{c������p�\_�o�X���-X��E��E�~�k|��D;އw�3�x��Vl�۟����^ȿ�t��/��o���迾������2=�?������f���`�O�w���<f|�߁�a<fK���$�{Q��>=Z�U�O���ρ��.L�ힽwLx)��hiOɞu}By��R��wj�N��~�����7��\��w���q⎵��/�>��?�������yџ���?_�c?�TI���Ʒ/_�C�~�s�U�~��k���!|���ތ����{����[`<T�u_����<e~��O�������Է���>��_i</��9��c�������"����8���K.�Q/~�㳵R_�^�.x]��GwM7X���O	�Kl�����~�e�;�O�3wEyǟ�9�K�x<|��މ�������s�o�sv�+��c����\��2�����K���	g��@σя/�D�ߣ���?&��V;|2��ݿZ%?�)���5y����o$��v@�g�;���|<�d+�7���G��른�wM�d����g?M�3���(��������=�/���c���菧����x��OD�^�Tؕ�A&�&o,$�~��������-��_��_��GN �~�����l������w����/�"N������Jڢߗ��k�'����'u�������%Ы_D}���ު�k�ޟ�P^��'�������Y����G��w!r��������c^^����?�7���Q>�>��OI����
������� ����1�>�?�^������~�/��c|�E���4x��~�I~ʛ��|��t�O�6{��~Q6�?���s/(Ux�����Oy05X��n�����_
��G}��t�˯=zF��_���uj���Hwϻ1��H��{gc��e�g{��;�?-{����S����V��O�8}7�~�5��;�����)�О���ϋ��V���/��-1�'\_�=�;�1#�	�D_�Lc��?d0ϋ�'\����w�__ӟ�x ��/rd�yZ����?�a����Ѿ���xƃ�ֳ>�Ş�^��'ȟ�#�C}��k����l�>]�}��������ěQ=z�F�����TK?�=����%��]�?�j��-�7A�x7;���5��Q��������iϔ���I�_��5��>Y�����?��؁�&1^?�!y~��t�K����I��i��3KV};�ݗ��S�;#�ZgM��e�3���z���ң��X@���w�����|r�����x��Nm�P�z:������N��?��?���/k�W3�T�?�x"}��������ҥ�&���uN��v�p���n�G����pW���������]P�������1���#�E,�S��c�����������{9���*{ ����O���??��������8�4�\�S�r���O��~߿������/&~ہ_�6�����Fz������@�/e�%��KVb|</��}���ο)�|=��}'���E��,�9�/�#��I~����o�GG���ї�����hm����Z�^���vI�������s����4��O���g�����W����QK������ϙF�߲=��-d�������<�,���r?��#��P��L���V�S>q��>>y~@��}h3�y��Ϲ#�w��S#�7�s~��w���_I}�o�~�ˋ�V��<�b��`�o$��'Z��ik��_j
zR?� ��G���?��=~O���ާ�@�g���*��G�.�HO�����B�;t�m=�T�y~R�ʻ}���L���[�&�񋧣�m��g��~R�|���/c|����S�� ���=��o$=Z��,O}��8�5~>���R�'���5���s�J?//y���X�O��x��$����U�M�'��<�w��T���O�W��7܊��.��W��ѿ�>-⯼�},����׺�A��E����_�t�`�7}�`��?�ǐ�3�����<�`������<~|%���l�u��0ϻ��.��_����R���%>-�P���t������l���~���f�膉�[O�OJw�{�g<O��&ǢO����i>{<�G<_H�ٰx�e�x��-������G6߉m���ևο;#�_������k���ל�+1�_����ϴ��>޴ψ���11��F:����/ǋ����N�D�%�w!���xk��<�H�P�8>5��������EI�����o��%�;���k穲�j���(���ym�9����������Ek���=ڷ�_��8~���7�s�f�k�}!�������r=��k�� Og��?�џ��������t���
|7ԟ�G՟�����h��[�kw������A����ܟ��A�w���7ʛ�}&���ߜ�_�_k��a�?_m��>����zi��_���X�ߺ� ���D ���$=�����X��翼����V��`�7�����^I}���A��(�A{��Oc�o"�hom�q�D����������7��wu�������OW&�gy=�'�y�/��K��|��k>�/�/棗�G}�?��t���g���;i����֟������>��F<ޓ�l_�,�v}!]�����������I~o��}>�}�?��������"�I��?bhO��5y��]�>��/�y�勾踿���N�(�����'����w���<�<����������?�_�j/f�E+	�H�[���J}\�{<���_�����l`���?ѧ�I��?�o�����}���K��$���|�����_��3>L�p������<[�y������'�����������K^�b5]��w��M����&o�_�_��%�S��|oA��d����=��٘���o��}ַ	�ג���P�d�#Z������w������R�_�>�O����c�<�ן��u����������}f4���}���������g�i����Y{��EI�����/����V����P����k}(�;��vM�N����~���-�(ۧ>�������d鏣=�7��W��)�����%�/m��a�ϻ�x7�^;�~��E���5�-�O�����p��~Z|��K���������w��ǧv���w��K1�^��)�-���#�-i��_֏����
��|i?s=M{{���0��'O���.�]����O������y�>�~c��Q�Oy���2�:�۹�}���L~�}u��1Hw��F�?��P������g�E�_H��z����1\O�<�x�?*,�����j�~Hw�f|��~�����t����[�����.]���O�����=��'���w�s���r~������;�=�4����"��i�O��}&���'��{�������~��<�l1�/5y��p\�<�T�!��KONڧ�Rg+/�?�����c���:�kO�]�����/����c�5�nO�ֿ�ϝJuG:�5|?��#���i-�H���C�_>���'~Os�������J��\�/�y�b�.�<����S�'?'�/����o)���#�OwO(�?�t�h��j�����D�j�ׇGb���3���~�ߟ����P�a7���q��b;wnO��������pm~�xYڽ�^����b{���4������'����������m��>�����ӻ�,*ೖ.޻�;~��coL���We�Q��=�4r}��t�Fk�/������Y�y�=џo���_�|��=��Ϲ��K%��;���35w��W����>��w|Z��Ǚ[{��3K>���ǧ�9�X��#s__�f!��i�|����ǋ�ϫ��9�w�,�����$�_���7��a���5�}_`�β�~�\e�_}��g�O��a�*�oZK�}��_c��kf<����Q�'��_���C���G�W�:�E���~��o���>����,Y|�B|�߭�;;����hϟ�gM�<�������I��9'���=������飵�M���z��t1���/}_x�����R��O~�=X�������H٪�{l�W�����xM���د��Ģ��i<]�t�d��K_���}џ�ע�Jҿ)��,7&��?�4�����������墼��wC�u�[�M��~�㣱�<r~������(��C�"��yޟ����DO?������bu��o�#����9?�/����e�8��O�e�/ܩ��f{�yt%)������L~�z�5>���������jk��O�L���p����3��/^�x3�����c��W�����|k�V�?��(�U��1>�58�ߍ�����r����y��E1��Z��c3�����q~?嗐���~���|����p���5������-\���8��ޭ�s8?I���bu�o;�R?/�������z{���S��җ�=�~������Ń�����w{�d��(��H���ӭxAң���}��_������\\���e��'K^����1����QY���;���u ?��+�E/�o�O�0�<�g-}��?ć����z��8}�O��O�;�k����c%��M3����V,�A�%o��e�O����j���G�=���}��4z���9��~_N~���@���E��qS����4�9�O�󋷎"=�?S��%K(����K~1~'��{s��q��b�]���|����;��Z��@yL��$����9�^��-�#�/a!��3Ӥ=���1��衷�'7F<\^I��}�E�-�����
<qz�Ѓ�C}����J��=1\�e������ѷ����暿���%�{~ٶ�^(���1��Ѩ��S0>���y�?��b8>^^�c��_}5�����җ��㭳����{y?b �����硽���ɻ�2����|V��\v�N��;��WV�V���Ƕ����d�3����kS�[����驾��Ǌ�|�>���B�7���_��3��F/�w{:���t��*������k�a:���#�K��s{��P�� �g�ŕf����J�V-]��G�>/�����)?I�mf�h�����_}|=���OW��]��Y~����Y�<���?����?�W|_���K�}�3�?�k�y�?������ ��	�~^]�u(��Ү~��^�+��|:��w�/[���k{����K��x�Ǳ����y:՗��[�:�?�����җ"�������OY������]s�o�w�-C���O��ק��7�����C� ]���߆������E��z��y1����6���<o�� ��@�2[S�����v���J��ɶ�,}��n��x��>1�7�U�>)O���o���_C�K��.�q|Z�5ɚ���mE>��6Kk��O�KO濡|�>��'�^W���Iy�g۲g��p~z�7�P?s�C{�1���b�g�A�)��*��ey��2x+���p{I�%�҉?���#[оt�GAo��X��i��l��O%=Z0ϻ�~�����oD<��m�.?���Kx'�a}/)�?)s���0^`����qy�Z~�7X�������%"���D����m����_���cª��=��w�W�*|�i���$\���R/>i�5�=ޒП�/Kve���x���?���R��>,�������y�������w�-�����9��~f����R]O���y��׎�]2�=��?֟�'޿�)��	9=���A�C�����f�����>����l�I��KOb|���~&�/�?у����������e��6з�<��i?6���5�}RR��vǇ�<@o�'�b����$���~�ۯ�>^-����t���?��6�W�ϝ�$kxރ�r�}>i��{+q��5���~���_�M����O.���]���1\�;��<��Kv�������P������d��ޞ�������������=?��nO_��>��G�ъ?��z�)�'�����1����yy�/yv=����OB}>��ѿ�I�#r�������Wx��o���b}�[>�a��%ܟ)ٔ�w��2~��q��+����F_߉�ܿw�\'��{�)���D��;އDz����������k~�}����G�?_Pr�zvE�,ނ�\���`��j�I}>�S�d�Z[�|#�������>5��eg�Qs��]�{K�<_�~|����%����	���,]���iW"�/���XK�]��=+|���COF����׿�'_��G��y���������%�z��C~��}���/�_��#�/�{�tңe/L�X������</[�7�o���ͅ��H���`�w�h�g�)��xx�׊7?���<�xh�]����\A���~�t�J2��\�|>E���E�����?���i��k��	ʷ��OM�#s�Z;��&����/[�/�}>��/��П�L�M�׳�2�����׏��x^��u�￩=�߲�|}>E~���|�Gi�_H/�G6����%޿�����5��� ;�������>o�Q�q<"��A��y�Оd������X{K�C~��/�m��ὀO��>?9�_�~����o�ϭ�*��ִ�=����?|o%�/�Ϸ&�q?��*yy�����x��+I:�{)��p�ok�T��f�G�����/��'v{����G����}_A�?���������e��}�����i�߃�=������������b�ukI$������zW��q�vE�k��߲)���<�ݲ�|?��,��3�h���B�Z���8|y��k����?5{�a�%?l�R߫XFy�se����G������j��#���w�>o�v��������+��������W�F�������	}k�k:�7M�w1<��9�.�q|X��诧�+�;�i���y�b!|�˖���ӟ���R��S�o�#3xg�Ǧ|��D�4�ˋ7����G{Y�����{����c����~ ��w�$���g����
��陭����d���nɾ���kѷ'4?]_����ϓt�祠�Z�?��i����ˑ�\Y���}ڿK����}�_��"?e�Y���s?:�w����s~z~����ګ��������5����+^��>�{D�ӯe��~�����_����GE���WG�~(���,���i�ރ�����y��{l>~��7�8=Z��~f�V|�q��߸�)\�&��|��s��k�?���_�I�����<��z���4X}��4��E}>�k�o�o8�{�5_���?�	�%�]�jn����%]r��7����w�+]���W@{����c�?�o��oF�Z�l�H~��������ѯ��|�~�{�����|�~�����޿S�_x���'��r{Cs��ik�����f���#�����?]��;��HY�z������S^����#���?5>��9)r�x��;��,��巾n
�O���&ȟ�7y ���]k���~����SI�^��Gy���)��6��W����*M��sv����,Z|!)?����i�?���0����U������k�ɾz`�>�;R~���d����d��7�{�WMP����Ž�/�x߃b�ݟ/^��J�O�Ws������ד�?�$���տ�t�S����t1���[��Ny����A����`��g��?�����?�x���\���q�9���#x�)8b��7��;�|?�������^��z߭�w������|�{GE�u�f�*ʳ��m�� �g���G~��h��Wu����O��ҹ�ݷW�w�p�i/d��������B���&c�i���w ��A�Y�9�'\�A|f������ħ���.k���Gȏ���Ũ���|���\s1�i\���N�C��W=��� )�������/���"�g��"�����j������u�Ky���w��_������./[�){�o�����[P�'[k~���}$���/���u�]�Iv'�i���y/�������58��&,��K���W���Z���4�>^�o��/�'�9���_m�q|(��;Q���G{���q<3yX��;����x�C�ߊ/g�����_������i�o��P~ ^�+k����2�ݕ����X��WƯ�on�*����:��9��]�=nJ^�y�	�[/��i������P�/�=�'��z������W@�?�y5���Wl�M~�j��ŗa/�~%�/��Z�.�p?[?i�y����'Lg{�>}^8V���[5X���u�箵��Su�� �sv��������`Ot?R���K��1�w\/�����������<��ά?����c|&�9��7EN��^mٛ�_���C��x�V{�y��O�/k�}}��1ヲ�'���ޔ��λ����8��?�i�7;�_�{��t�)�Gz��a{\ߪ�7&�`�'=��["_O�/����(��w?OKW�/���4�<�3��>�N���'�c���x-���x����>?�oD�_D;�O����+��SK���C{0;ϡ�����^��ע�f�6ƿC}G��|�~�����w�ɤ��x����ߚ$����}(��zej������<����r$����ֺ�ao���}�'@zp~�p<i���_��h.�q�x���s���6�~��f�{Oe<�?�e��Q���?�/�E���^��z���IY+l~p��?�e}E_v!���DSDn/p?Nk����~dM~.�8��^v�!����/���m�a<�$I�>q������������O������cƣ�?ꟈ�㣲�����x��>N�m�~W��x�[E}�~��[Bz�>y�/�su�NXߵ�]�r~!�y����X��O�wN�'aj���?>5~n�G�7߯��ז��|>�.�?�����_J>���{A���3�����L�Z��I}��u�����8��1<��菇���IV�����[�������~"�ò�?`�0�/]����h�;�������^�?�����1n-?�_��V��?���]��se%���5_<^Lc����^����r�n�Оr|�w���S��'��>k�����c}�o���-]���W�r�%���=um~��,~H�|��5�^��}�z?��k>�|)�f���,oZ����_���@{�|���pW���ͨ/�`��s@m�D�&�Tm��S��֒������B&1No��A�[��j�����'���㝹���7���?��)-����B|���u�X�&�oF�1���Q���U���#��ȷ���;�_�߼�2@/������?�M<�H����/�w�G�6X��I�>��Ux_���w�`�*�'{}������B:ק<����5��6�߿�x�5�gR>���V���s�v��>�q���9��^&?�s����3�����z}�Ħ�.�~��_ےw���;�������bD___��3��I��ߗ=�F~�W��mB��~l$�-���"����5WzS�H�|�9=�{�J�	�Z<\�������j��#�d��1�s}��S{���G��[��#8k��e����>�Η̟��5��a��gho���>�����C����#���ob~�}H��y����� �}	��ߍ���\��x��S_�����#קZ���R��,���A���B�����b�C�7������~��=a��F���f<ϐ���>��;��G{/�^����.Y���gS���y�͵�@��C}��1�������e8>���{l����.���We�{�u����Ψ��O����+�?�g�w+�L�г6N�m��W�����`����xfO��b�׽�y=��������۵��N��gR?����$K��� ]�����`�;����w��/�y����ί���f?�_���~�"�o��1~�"�G'���j������菏ǟ�W3y�����{������2}������D�n�<��ޞ�+���ć�|�;�ђ'���>������|=��+����m������~ˀ]^q?��}T���>��*�c��?��L����������}wvW�A�#!����Jd/�V"�f�d�@��9� 26	08`0��6��lcc>�8����8���:]g���/����w�T�{������N��������<ϡ}��0+����j��ѿH`���kI~�Ͳ���k�/iof�7�k�?G��A��L���u���{Ԟ��֋���$��p>���g�yǋ0��ӟ{����y<}���?�������^����q��./D�/���#�ۏ�חGE_ޓ���{�h��e˺�`�k��Y�8a�����
�g��c�����Y3��v��7�1������/N���j�.�]k0��'�����B}����?��j��Ǣ��,z��s��k�l��
~���I����'�y�ڧG�ߝ������no�y(�菗�|���+�sz��gv�|0��O�JV��I���_qn���I	�� ��׶��mo?���#�����O?��|�������"�O;0��k.kM��b�>dƿ�G%�������Ҳ�q��|�:�	����E����|����ݠ��W^������a{�_�?��O����*���zy{�o�A����p��1�o��5���[b|��|�>����J}ܟp?����5�7���O<��~޵��?�G�L������d<�i���|��wS�}���v^F�q}��S�u���9P�+;��������>zz��	�Z���O���/���ˌZ}�o*�bp��Î��ܟH��R���>�7��$��?iK����|��Z�y���ry��g���[b�~�������t����o5Xi|O��3ӷ(�g2k����]Y?������Ǯ��[�A�οA/������?�5ש�g�Mz����}�p�~���]�GZ��H?��=Jϵ���ݧV<��&����]�I�;]���n�����0�x��}��f���\��^^��6�¿={�KyG��ן�h�f����R���{yR~S���<��=�}���0���SY�]�/�_*{���1�'M{Ϗ�������W���ϼ|O�L�Tp���-����2>FT���g�rl�
W��<�TA{���J��35�m�?b8����%�������v�ħ��;�}͍;���EX��x-7"6�O�?lOm��Mg�~����~��[`��o����W��.9�k�wy�W��c=��Ӈ�Gb�>P�G_�?ċ��;����g�x�8��ڝ姽��%k'��<�������u}uo�'�W� ������-(_i������_C�N��ӟ��2?�'��C���pYO�e{5����O��J��D�C�=}-��K����	z���݋�t��_i%~ԗ�ޠc|e�����1<�s{�����(�O�����x3�D�<~����Eƻn��?�����>�I/�O,��ş���O�~H��V���%fp뼐��/��������9����_B��	�d�d�/,^9��'[�G���ܤ�ҳ���L��(��d#���km8
�xy��퉡���/Y����G��~���n���,���^��<��g<C�'���V��`��?&�]��}+O_Fz��5��/f�j�����3�V��뫼�6��X}C�A|'1>��'Dߓ	}j��?������d�u(�p�.z�z��x��Cy{k��W_ꃵx;�=��5{�����}�_�G�K��/�l��B������gQ���m��ڑEo�����ړ����Ẓ��ߡF��[��_B{wM����0^��3���?���4�܏�~d���'����/y����?���#����<�0�����ӗ�5����&(���5����/p��^��S��������8�����Z��}lR_�p~g�e�׫�h��^�^k����񟂾��g����x���Ȏn'�{:��B���2��|����n�8;�����؞��|�^��z�>�_�Gc�I�����	����̛�3�g5y���/�P_��9�k���{:߷/<������\O7���5b(oH���,_�b��Hj�P����l.�z�ُ��}���ןfe&��`�s˞�������O������I%���?�oPY�?3A}<&�>�hwe�~�� }i�ůpXe�^��]>�����-���]ͭ������H����_>��0�ѷO�~�����S"o��9���������~��~���U���+���-}8bh�uzJW�&�U�7���6�c�_�3���/&����z��O�q|k뗟7
�,ޛ����;��3x����E���i�1��A�����^��G���G�u���[���1>�)������|�T�/:=.��y�c%��������}�e����	��������1��?��E}렷�'z��!y�L����j��|�Xs�(O����������Ŀ������W�W����~���'����ħ���O/ �q����ϵ���|��mͿ���~~#?��t���ş�ߩ�ۛ��^E�>�i�
���ڼ���їg����~������ZҲ�f������R?}R��v�Gd{��%>�������.�Զ���w�߯���l���uy����/��q���[�M{
�g���+��;/�}�f�����B�g��2�{{Ǣo�����O��>�y���y.��пeЋ�i||~��O��7?��xp������>��~��6�|�>��k��ߟX���A����x�k��Ǩ��_!�+�}��i��5���7i�3�zo���r<Z��N��L}��X�o���/&I��[O�[�������s�_��Yｽ�+��ch�ҷ������(O{����=��\�����.�G���}@�ϡ��w��x~M����|�y�ӳ��+y��9��~y�T�lo9���?�g:��ٗ�+n/yGi���r�����w��2�vʻ=��Kɯ�7�/�������?��?��,~_�v_��u����o����W����"�!�6(�}�H��\�`}��K���+d�Ʒ����ϣ�����}������kz8��Y5��M���s�h��ו&~��������h����Cڋ��[lOg%Y|ˍ��]���� �u�"zg�LI��Ɩ�Z?�'���#[�_�������5�ܿ����/^��}L�ty?�����ыx"I����xߵ�_�>���l��x�~?�?w�����U��֟�h���e燒�7$�m�_�s�]��^A�ߋlٗk��-��Qp�O�(�o��)-�j��+��J�_D:�K~�,��9i��'=U�q��{���K��	�;b>u���76�]F��b~��ſ,���$���>Էy�/��z��sҀ�?�������<�ߔ�����?����$�-�/��e�j�W�?k�8?�ߏK�����IzM^�#�gud��Χf}p�f�i�g���t��.o,�O"}j����%�>�4�����?=V>��q���Q��O��|�����9�G�x`�z���_�G����x�����g�R�� �M OQ�������)�Ə��g��O<���5W�����.��I����x�u����7�s�����a���P���:�����,[������}�[�P���Ϗ�>���ӯ�O��j��G����_���}�@����_����K��-���ۗ�vy�9����g�ںu�޺#[�m�����������,���>�ߓ�S�-?��X�y��'ϋ�?������P�G }��W�ܴ7p<h�wy��-џ�|O����C�KWs|+���/��������[�)��?b�=��O�%k�7��3ۢ/��}����?ύ
��$=@���'�ǲ�ڌg��;R�=I��r�N�9�������x���l廒���}""�_�1��g�<��髹������,~8�����S�7����˗�|���y�:ks�������ӈ��uj���;�Kv?T�c��_�z��Q��㽀t������o�`�
�o�����~��,D|��?�_�/j��y_'������sg�����������_-����|k��?����x>����I��������o�]�~F���/h|=���@�X��'wg�i��gs"���=���may���Y3ㇲvn���K���1���Cy��G����uN�i���j���K=>�h�b������\��H�tQ������_���/+��D����#�\�^A���/ܷ>�>��ْħ����O
��P�~4�����̲7��~�o��?��S�/�њ����������/�����`�M�A�\Ϧ���on6gf��bO����_���1�A�/��.��&�/��oh������d��j��K[�H��w�#��,[���|I�
�'h��N���0�t�%�L������_Q�O����Y�
����}����!�O����k�u�_}�*I�ږٟp�|��99~��u4��שH��6X����������]f?>X�߆��}��ӳ��c�������O{�w�=�������)��=V�Ny���,�;I�o�������C�g��ǯ�K/��p��u����T���y�k|����i�z���J����g�}����-nO��O�YN/�C�^XP0����{��G�O��������E�i�`��yI����tڇE�,����?��� ?������{x���.oǩ����������}��K����8�f<��~��4ӯ�/��O�_�^�t'�[jٗ<]����g����>��vʏ��h�'�_��ɤ~ڗD�_5X���W��Z���������H������)�U�y�F�e�꾪AO�cV�����6���\��|�^+����puR�/�О�����|�t���v�MB_�����<;7)/^XA:χn�t���r���k��=��_�~�}�������O��/G�x���L�g{��_<��ݟT�ř���w�����k���`Χ�1�����Q�/r��������syD|��l��\?���>����������0�Ut��2�g�,�˥����9�Ї�(�y�A��c�}��|�G���+k���A��x����!��}}xA�L�﫹u���ϟH��g��J��n�>����{�wͳ�m�������kj�ON�?�����_�J��~��'1<��|��Z�z;���^�Ok�/,��� ��T{��.�=��x����i�������P��%ߕ�>��R������3��_���Q���O��Yi�t��?u�q�K_�����xd0�cS_�	������pq�V��yw?Ǉ�;�-�'��A�R}~�Bzq>�`�_��5y����3{�K�9?H�|&O�Cy���`��3������?!->G�|v_��$�x��x��?�7�/�?�O�[i����+����H�|��WRKv�<���>�5�n�<=r�h�p�B�-v���y�]�#�į\��8�tޛ�Ǐ�k//�=��#_&�g9)��M�����q���`~�gZ�?ף�����YK���'���+��{R���}q���t��&�����'���K��k�>���K-���w�?�@��o�~����r�Fy��M�=3~||3��� ��\|]���`{�Ǚ��������k��&1�>�Q���p�����<8�z��G���+��|����Qo�F_��c{�O�<���9��xj��I�Ny��S���?��?]>.o4�]~R>�_��ѿ�־���+�`��b�?;_��z��u��������N�|�<��}�=����S�~�Q�y��|���_&�W��W�.o$K�d��/_�۾5�㗭�<�ٿ��>���+Kx<9���,}S�ғ��2��z��'��u{���d�>]�.d�-��ݑ����v��X?����H����/��Hҍm<N�M��f����+���Lu��xo���}�F�e�r�ŧ�_�~������c�OK�����nS>p��Z�V��l=���O�_����Q�3�����D����&?��۷[���|n�t��������G��u�oN҉׋'��Ǔ�}����w>���~&�'��tEw����h�����z���������Q���H�2~��w ��{��zK~^��'~ۑ.~:f����㑿C�k%z�|�uX���~�?ϧ�����h�yw�߫�����Ao~���_������4�畔7^_�������O�{����#{����kS���tKvd�Ư���/���)�}}X���A�|�����������']���.��ѿ����c	�-��?�	�����y�HW�|����W/��>��>ާۇ�į�����v~���6�����o������x�I?��~�5���%��/���j�z~�^��罒?Y|�C��C�z�ڲ?�x���2������gmf�K{�W<���N�������HY��S��~�$�9�?���s��ϕ����߷��?E�;��t��w}��1��O}��������MFOƯ��P�����쿭�M�����Y��2���1ܯe��+��%�C\��-1<c|4��
ڣ<9��)Ǘ�g5��ў��!���>�O�����B���+��6���s���ߵWX���-]��Cz��7�^G���F�w���L�H^��t�vo��I�⧯�7�n/���;=)_�^@?o�-�g��������+�}BR���E�w�w5���O��5�e{9��?�z��\��Bz�����G�t/���-p��E$��Z���3���U���>����dׇz��Q�������|o��#~�����������Q� ��w��ܾ#y�Є%��O�%�=~Nk|X����3^��'[���T�{�C�O6?�u����Ͽ����E㷖�g�c㭱����/��K1����<�?�����˽�/'��.ߎ�z�>=�sʇ��������V�[R_R{�_�X��5%�]��}e������>��{�=Z��Jg�����6"�G������e&_��h��}0�痢�G��!��/G����]���z����������1�q��
���O�����z���]�������".vD_�C�����'����y��/�w����>�������r����>k�����C|���p���-{���_ԗL�n񫾷M���C�}�M �g���;��I:��~%Zf���~������j�3���R������߷������9�7kk,�h��}�w?�a��z��O���C���˞�#I���l�������t�P�IEǗ���?l�6>�?ϻ�?u�X����|�n���/z�N���"���L꣼�٫<]?ޟw~.S��_���:`��۾_���[�/O�1�w�7�/��b��_1Xk�������?��7��#�N���[�rz���9��o��p<wD��*�Swc������������-��Y������W�|���Yc����ɦ�w���/ᖽ/4��|�ڋ��9\hًV���/x���h&��~�>������$=����`�������!����(U8?����~��{}��1��m��x���2Xcw^��7*�0����h_���P���7���$|]>*��n�EK���m��<���H6x|6у�����VIz�P��$��?��4-��`<�x��F�_�"�OT�WG}���0��?8�)�x�7�~.\W������\?���)|��Ds��if�,��6Է-����1�/��_���a��L?g؞~��(��w�I�u���t����x+������e�>j��&�s=���7�c(��~ɿc���P?$�-���ۘ^�ߒ�7�"��|}=���������3y�a
z���3���;���6���p���]�ų�E��n��z�r��&n� ?j~�����?�����OXm�����]���O����-!�6?�����x��Rb�̟��/�칔���������2X�\�_��4u6c�7�J��]�~������������q��>"�U���(=�$�O@�%�������m��F{<_9�лf�px�+yy���tM���o�#=�^m����r޾t�?H�G�e���gv��v�_Q��W�����~<���B����_��?��J��8my���N�����A�_c��F���|�5���#q��[��<���h���q��'�hO ��? ������O�����o�/���?�Og�O{�3/(�w�?�s����ҧ�w&��k������N��.$��I�#�4�/���~�o��?����?{��ۃ�M�?�3� �߅�z���خ_��ek|����"��ׇ$������s��ћ�����a:����3���}�=�Ok�ǒ�Z��5|������I}�������1����Z�~�`�ށ��>͕?O�W}o4�ߖ�˱$��s"�n�<�����;��9�뻼�ܝ��g%����˷��#����op>�	8{_��{+������W���g}��F�C�_��y!����Z��<ߢ����m1��h���3���e��T���H�	�o�k��l����d�a��Kl��5���]��Ygc6��џ��sG�����/a���(Ɵ��{M�b�h?l����|v�y��~�8����V]~^ ں=p7�E���P^��g�A������|o�'�;���D���C���=��[�J�'���_�Eo�����&�G֣O���*�鿁�)}W�ӫƿV~k���+�V��P���x��Ogs��V������.?�)��?�x���\ߪ�{���{D��u�����:����,��W��s|\^k<?��Ώ�G�m���.�d��9�i��y�k�t�[�B��r�P_sy����&Y�o��e����<o���^1��c�27:����5xO�������L�/��ߑ�K��}�C�"_�Z� ���m}"����������op|Z�K��j�Ǜ��L�i>�~W��O�<�e�����$����R�H��R�z ����S���Ү���������������Q{��ז�F}-��h��ܖ��X��:���y��ϟ�%�2�G�[����Z�0��5}��u����w���N�����7eIڛ��j=f�M/��r~{�~0��ᡠ�J�����B~�����;����"����c��t&�+x�<b���������_�~�b��d�P�a��˫��/�j.����)s�s��������|�<���菷d����*���cO��O�}���]_&>������������,��0�o`>)����q�~;��N�y��`}3���	����|M>��!������F{:맽s���]�|����+CyI{�����k�]_Q_�g��I|j�;?�n�������_}i�����������޷�������e�ߙ��7��>�����+���v��|ݕ�K�6����k���/Y���'������Z��o��#����A?�7��{���m�/tE��d����z�^���`�g���Iv�X�q����Ѳ�_�$�|Do�Y�oA���j�[߭��C~���Y�����O�޹+r~/uu�h�h��[�?�o��I^z�S}/Fy��XNҹ?�>H~��9��O�<��ū�{�܈��9)і���{+��t��=^�֞�,~r�����="�{>�'|���o����&�<�|���r�;�~��~v��������'a��)��E�V< ⷻ��l�k���`��}h�z�`��{���+������/�G�t8���OoT޽�|��-���&׿[��L���{���>�=
��{r��0�[�,�=�>^���>�T�%�����߳W�ܟ��yE-|�u|/�����g#���Ȳ^�?�r<��0��]�o>�W����9�g����J��������ś-�����aI{�(�u��Z+����]�Wb�����A�f�~�?���ˠW͟��]�x�����7�+%���^����$�����/]�.IzD���.Z���'�����~�s���x�5z��\/}<�7�5�g<1������	��֏�̷�������C:��>�����i��l>�/O }�/���K���,�\�ԷO\���5�c����nľJ~�ҝ�ܯy�=�`�'�>�Z�y|
�'f�\?�����%����[�O�����ǁ�(�����������[0㻒������7X��Ο�ҵ_�,�������|?Ky���9�����g�����I�E�tگ�3Ho�'�g�z�ɣ��|v�����<��wD:���~X���%�l��._՞�P��|�^�sN��7$��,������%|h/�t�O�^)^��s��}�\¼OC|�/�}؈\�p�_�w�'�����~�([����+�.���C{���9_���^�G��_Z+ܞ�����F���Ų����o_��zO���Ѿ9����x�?��#��E���������h�/z}5��z��s���8��/�������W��J�uw�7@�l��-��{��ی�N��<߫��E����V����s{�4����f�n5z{�����颅���|�o��{�Z<�l=S~?��<���x��b�=>���}��?�R�G�pv�_{?��~ߊ�(��U�O���{��??��@��9�ٲ�i>�>���}3�����z�~���������IK���o����D���_��O�>���}��%O������f����b�?��j��!���%��'��W =������~D��6�[m���y��e_s~$�[����QI�J��W- ��/1�g�>�g�:a�@���o#ߓ�wzɟ����_��I{����C�g���g��_L��_�k�ҿ-���y�&��_�^Z������������?ǻ���Z����诧-�,���Gy��]B{���������O�~��'O)��b��.?D����׋�۟�����!{�d����J�!I�< =�>��X��Q5h�o;���&1�o��� g��"��[���t�/?]���n//����9��������gwE:���4�!�?о�^\�2�)��/��N��gK�O��e|;?��\<b0�K�_?��~ ����o���^k/�B�������Q�k�_�o��h_��5����'�>ޤ'��c�Y�K΋O�=3���s�}�~���������>J����2���R�O�غ>���ό?K�(��yj�	��ݾ���;�O~h�C�M�K~=6I��ڬ�٥�O�S��#�?V�,���Sx�CX���/��=&�Ek_ߟ[>_N����t�Q�[����S��2��x������Z���j��o�=bO������|!�����;������A�%�i��	_��U�/���ӕ~�҉2�}�QZK��{3���:���'�_��χ�����]S������`��G~�~���1�{t���Mų��͌��� �K�q|���3����_Z�~�O��%�?S���;������=��Q�g�"}���uM����#]��9���7��Y�����������2��ů���`~�+�OVc���s~Ȗ��)i��z �g��]����+d�,G���d��g3����{*�����n�+�Mc|��O�>p[�_N�K��Uk_v��0�s����1X��~�R_�Wh>�xL-߬�]I{5zr=��4��%����s�?-��?8��� �11^?Ǘ�������3��>={w�,Я|o��o=���\W��b=��B-�����콴wd��u�o_?��p�ވ�}?E�T݇P�}b���Sݾ_��A��i�k3ސӣF��q|5��=��mzg����zC{���V�9�G��*��Iy޷"}�J~�����wE}�?j��z�����ӑ�P�_s�����w�ѻu7�/;�����t�%�k�H~!��D:�;���h��֏��-�/���1*���C����������e�ӭ,�}����碼����>�^|x�3�������9^�{laQ��Ez,������ۛ�/�;�ȿ��燖���)��3{����nV����H��R���?2���k��?�F�l|8)����� ӿg���3+�;����|���;��/W����G��Q��5����G{1��k����(/|��u~Y�~<�Ѓ��"�>�������?��_�j�a�b��7���y��g�88_��߿���^�x�	\���-}����K�8	�/��c���#�N&�1���Y�2����Il����+ȯ��b�~�e\~,��K�/Z��*�&�ò�{-yJ��?��??��|��lco�^�X���Ҳ�V�O��Ӿ��],k���/����o���W}��n�-�W��?ZD��D��~N���c�������,!���E�~[t���׿��$�����_���1�OQ�?{��������O��By��p�����'|o#"����v��B|~�x<��ǋ���%�W����D���v��^n�l�oC��|^����(���y���%�<~qm���\��ן��,|����O��q��~�F��-�MyH�о�����*=���U����������x��o9��?����߇�ޜ����xe5Ig{������Ь�?���x�����g���M���x�� �����S���g���m0�1�'	7�������Ҿ�{i&�����H_�G�c�~���^I�mկ_vߘ�������b<bއ�����*E~�e�5�ok?S��_xfA�,����G��_RcG{��Iy���N���1����7*���2}a6����3������?�z����~X�_��3����~·������q����ϧ������ڳ�O�Ύ��~��6����Δ���>;����s?�����]j�Ǝ��L���Q�}=��`�1�]h����<oT_hO��J��οg}���?�z��?魵����e�	��^���	��#O���)I������z��a��{Q~0�����|�}�F�ߌ?#��}������`���e$��T�+�Ok-���3b����&��S\nD>�|�~�`�/|??/}���C��;'�EO�w���>1��mv�_Y;�����w'�������_����䛾����{���$���_ӏy>�����'��e�sgu8=��؞��/���yU�/���ߗ�k�˵	�������O���V\~�^��w�뛼�,!��t�W���$�\�\oy�����/&�Y�9��,F_>���w��em�V�z���G��,^�?�?�����}�)�ߌ�V�?;�Q��|C��M���K�r�Ls��Cu;?�+�gc��- ^K���sd���R��O���A��}����[���U=�Z���z<���uk�C�e��<��������V���������xY����s��h-���|=}�G��n/�������~_�`���5�g������2��tK�o%=��-'k��W���l�[���_{uυ("�I�����E�@������/�^}�>��}��{Ao��S~i���l/�����h��}=��w�=�G�g��f��C�=�Q��?�ҍ������6�3�a&S����^{�y1��;?썾����?��T���,���b���Z�ϛH�Z<Yί����Iy�B||d�xP��#�r���J�n�Q����K;������ǃ�����ۣ���E�^vF��mm��ڟ~�lu���_Wc�?�����?�����Oy%�}>ʳ��+s䯽��5�
�I��u��U�V��>��ԟ�^�s}���ǿ�/���k�_��K�8Ioɏ��������<?��=o�����}�_i�;P��R����]����o����/G<�W��7r~���lo���F|�zj��K�߇R�[-����{|��W��7����V<�����<��=~)��.y��i�'�O���P5|=}�oW>�� ��7�������3�B�s'���|�����/�# �����?����g�p�y'��3���y��۸�����[��~�V8^��yI���t�����?�c��G����^���g9�v����o�_m%)_�w8F�Ӕ�����Q?ۗoԯ&�_J�,�~Z��9�r(��n���������f|�9�W�W<o���x���6��N{�F���!��>R�OH����n𾯍A/��� }���ٿٿ?O�zoC:�_�ϱ9��'~t��|x���D�����\��l��%�?��2�s1���Z�㝐�t���a8��Y����6ʖۣ~�r|E?��ތ���WY��Ӿ���؟��8}X���
?���y�g��՟�_����ҕ��<����u�����|���?P>Ѿ�����q�/��S�t��������}��<W���[��q�Ǟ)��/����$��\[�������0<fs��C\�gc2V^i��mF}�?O�ZIm�_��1��3۴���?���S���9��[X��I}���f	���b|/��2\�h����/3X���l����5{ߧ���Mn.E�_Re%��3"�_X�e%˧���/y��o�\З���(����������.O��`�"���Wv��x���3>bk�`����G�>�����b{5�mfY�����X��~��������3�Y� �|/��)��>�Gc�f�懟W���*燻����_��������:�)�ch�d{�������g\j�����E��<�y�����+�_??����+��),�������ᡀ�P�{<ɍ�� �5��������:�����;����1]���|˾S��]H/����{ ���ú�����K������T��l��
ڳ��>�}��6gg�@�o���\>�?.���:?�n�U\�]���#)������������������F�����h��G��~������G����O�xz��u���}'����$�'�'H��4���(��7��P���\Y�����1<?�>��7�S{s_O��u~��ו��N�1�g�����+e����ڛ����˾��_�����K�y��2���.�S)��Y>^5���w�[�᤾���a��h/�?�~~��=�I�V�ȿ�?0�>�C��y	>�������7�ϻP���Ok���d�������}���
�g�axߕ�z��Z��C������{cY|a�ƼoI~ɖ��t���g�>=�����k���ج'���+��-'�k�Z��e���-*ܕ���wy!�F��ٯf4��*��m{�>ο��>�7OK�ُ��qzF���<��}��}���QP���=¢�{A?����E{	�A�'�e�o�75��X�_��)����������3y'\OίZ}��y:�k�ۻ��0��O�����/�#��0�T[�Л�5��'�l_�v{)֧�����V����P����l����j�[�[�~��]�O����x�MH��п��w���0��%�(��_8L���]�[���Z'I�����vx|��F�YϿ>Y~/E��_P����~�e�_wnԯ��������*���N�j�G��g�W�_��g�?����=�C�����t����Z��J����!2������������7�~�ƛ�7�_:?����g����0~��zd��'���f�G�,����������I���KI����s�~��'׋̾����_���_���kn��B�2Ǉ����@}rW�%p6?fs~������`��Ͽj��7���x�*�M(��w�x�=��35y����W_�4��B�>�<���;[o#���L�<�����c	~*K{q�o�?WG�D���=�׊7��|�t�����<3�/��_5�(��o�(����`���=!�h��6�����Cv���d��	��������W��^�v�g"~ޟ�/��h�l�ߛ��<�����A�>���; �f��C�oR�p>s~f�������/���E�M���[����5}�忑٧��2�Z}^^s����W�1��?����0��Om��>�W�+��4�D�}��e�ع?p��s������G~L�G��֙��bgO���>R~��c<h_����$�Ƈ�J�?v�QH�x?�}[�?�|��_���\t�C+��3N�_��wX������^1\/=?��E��,�t{3�߫
�k?��7<��{B*���^�L���O���`�7f8�`��c��������cb���
ҽ~��#���o�w	�7�w�[�~�7�d����?���G��\����ҥO���R��_dGg�/^z���F��G��Xkٻ��r����]���{ ���=���(b���=�񗯎�k��~�R���C��~��h������j�������	�_�ݵs�!�D��i5����C����46�����D<�=���[~]�_? z�^^���S�G~�g������ee[t�����鏪���Z^d�2�1�g���@~�����e<r��2��ǣ�<���I}<����O����>�O��|j�A�G��<����#u~r%�s~*�2q����z{"��%�A�f��e�A�^��&�T�O���}�G}T��W�c��������F�Y���|}�Y���?^�����}a���}a֦�������}�m��x��9�cm=p���|���6�?�m��-���V�0��ї�5y���$����'1���������#��p��E�|Om�����`�j��S����=����#��D��j��$w��xtK�;!��?�����������*��I	o�����_H���Ց�W��;$�G����ٜ˿}���c�Z�E��}��	߫t�l��p��}�Xt�1���x6����D�_9k>�>����o%���x�㽳�wF�|����_�u~�oC��W�]���(��O�ȿ��3�O��?��R���?~-{W�>(�ա=�GV�o�������W��3�'��{�S_}+��Z�2�K���xy�a�[m�>}��>b����?��7c�w�ל��3}��CX��v�O6�������ܿ��%��?��d�[��g4v~�~��o�<Lue��4�+[�������^d����I���B/��������L�s���'�^X>O}W|[�`j��Z���k��i��z���E��xk�L^�/�什��K��dR^��'�u�/���p��x(��(��?�ߪ��|_2 s��}���a޷��?{O��>3�������菇dϵ�wo���D����5�'�?�/��������]�����Lޒ��2^�C>�t��b���Ŀ���+����(_��x}E6t�o���4�_s���y^���p���g�xz��s���׭��n�~3�|}^��W{����\~�I�w ����H'|f�?s~y~ɋ���~J�L���Oc�޼��e8]�-��>���b����s�2$�_��y�J�~)���z5���Ϣ���<c��xv����}&�I����l�g�~��>�O+�P?�|��ն����T��ʻ|\��^1���>��� �σ?X�t~�k�_���O����/�S������s�>�#�.�6�e+pM�� ��n��G����k<$�w��4�|�_D���Wv������F��*�9^.h���6��~��?�?�K��k�?�|��gMx?��������)����WHo�7����d�	��~���������'�Ѹ=tf�[�����}�G��W�"~����]����~Z}w~�oa��������i�h�/�U���`��������K/M�o$������o�����#����I���O��z\��������{:��'~�&�7����?_/Ύ�>���y�sQ_k���K���1^�l���b<;��eK��1�������vz�x]��{��/����r��x0�Cm��o��\�{|*�j�ǅe������J��o�_����'Zx|[�����ɇ̾*]�SH��S���\�>��������5y��w$����֒�H���U��B����%�8�����%��K~��y^��K~g�o���>���?����Q�;ӯȏ���~F}�2)�x4�'�z����s�oߕ�;��x����9�����a���5�_���sc�{���]�2�����_�}���>�_{�����ҽ?�Y>���_����µ�w|�������߫��E�:�ͅ���R������_�{����rz����>�2�"�7ɖ.ο?�#}�?����-����|�?ff�}����/Y��(��-{���L?V�~�$��	�k��L��Yў�,������?�f��>�ǹ�J�ܹQ���>���/\?�G=���?Q >+���$�;q�Q[?'���o��S>�k�}�}(��Kk�e����.�~?O�����������d�3I����S��O�礿E�������㛊?���j��>�<��lw��Y��o�����,މ��$噟�@��D?;�s�����-���s�=!��0�����<�㵐���8�?s��,Y�����K���~ؽ�d��-��(���)~q~�����O&�G������|�r�����=���pp����E}��e��}������1��h��Iy��x��#���9�?�������%�Z�[0�K������*��0�s}Y���F��]���z���=�w��y��uWd��*�~���o������iOk�k�C����>��#r}��g����k�[������0�A��o�K�L_R^�Ϥ�?���'ԟyq�_�<^�E�}��=���x~�;��	���s�?��
��|?P^�:�g�aD���� �+���1���0�����ߚ�~ߒ��|���$}9�m��]�P����e�iL{[�>���;�o���|���ӿ��l��%�]��f��e���a^��诇?R������k��gړ,�������+҇�5����4�6x#�e��V��/����� �W��>^��"�g�}U�������a�oƳ�������'�w޿��z^��<��F�8�l�<O�}�m�gK������-�VM�s~R_{Q����믷�����x���Z�~��������P뗽y�O�M��?\d�x�_!�O<���F����3����ٶ�S&?�}���.������;��""�E����NED|l��xy�Sy]��������m��a�?/�/������H�~~򯡿6U��Ǖ"_�t����Tvj0�'�>~k��%���ӗ�}Ho�׋���Wn�W5x-��q~���r��Eҹߥ=6�/��R�[)/3zlF�i���h,x�����}@��s^���������3P��Y<,髫�˾��'��z����S-�p��������8�!�;�D�C����8޵����߈�ߨ���2}B�����'|0N�i�������ϗj�'Z�3zP����x���ˋ��矯�ۢ�����4�n�^�R�W@��Cg�C���� �9�i�����}���I�>��^_����o�<�1K��ڿ��{e�ދG��n�����?���p�Y��3)�ؚ�w�����I�l���|3bho��W���'����ߊz�K�o:��A{5���1�tV~6���������������繠�?g����{u�e�M��;���}��o�x5�O��ևc|�)�5_�}�_-]v�3b�^P޸~zUi���ۿq��o���5��L�e������6ӵ�?�N���O���cK�W���V�o%������Ǵ�5��u�_ xCypϤ|K��}�s|4�� �x �����G�c�hy>�g���q?C�8^�O�h�h����|R߯3X��.��f}�������Ʃ7�G�S�?wM�C���C{z�_���|���|l��ɾ���_���$Y���:?�����>??��[����wC���/)�C��/�G�:�D���{磯wkя/t�TA�d�!⿦�2�x�I:��Sgso@z6�HO�ֿ#��1No�f[��ɇ���K�?��O��l}��C���/�?��О���kҾKyi��,�D���3��K�̿�Cj�_ߧ��o�z��1���+1>~�s���c��ղ����g�F&�>^��x`���;��r�����ϭ���x�����}�����������wfs����(���=����)k�ΟK�����?�W��s��$+n�����W��W���2>�#�_���ɓ;�8����G?/��\����i�5ʓ~����w��w��෗,/G��#�_|2yCX��<-������Z��o����}�����a�wy����'3�`�������������ӿ��S���~�bp�~���}��Ƈ��[x�f���Y��}Es��q�u�������ۡ��������e�c_T>�@}����*E6ON�~�/Zސ�Wdw�)���|��$�P~q=���i�Q_x�s�`�'ʷ�G�{e������HɿjoR��E�i��/۟|�4��o�;㣬�<߻��Z�� }6�?�흻��>�$3x��ǳ��K��ӧ1��=�� +�=b���=�ofo���K}�|U���I����ů����>ْ����/���|I����G�緒�4�����w��B����ۡ�lO���V_}>��>}���X�Ǭ��iѿ�:_`����������D?�o�?���.�?�"}&Sf����2��\y���*����W<�?7��=�{�����W��j�����,�;��-�}�߽$g���_�Kv�s��3���I����ϵ�X�'|=X��}�������ze��')_��t��������ϙ}�&?����<�����hq�_�X�>�?����B���w1�G��?�������~���؏���������~�&�����./D��"?�8��M�|?��������G�"��<�"��{�y<5�[m|��"��%[�ò�t'�?���p�{J�Gb����`��xi/ꧾ�������F}�����秿�-��w�����u~�������^&�E{�ߊ�����Ӟ��~����-X��_(��_Y��m��L���~ޯ��L}!;�⎿*����D���|����x1����{y��`RD����<���|?��D�?/�; |��F�4��d��H��ޚ��k���S_���������/�����������t}����%��_-�a��Ϡ=��Ώ?��ؑ�g�
����W������w�a|
گ��#Pڗ:���h����v�?f��m���7�~|�W���g��kѷGN"�H�����`�z�?�Ɛ��G�e���V�������GPߤQ����w��ʎ�g�w��|r���[�[kԟ�ok?�-%���h�����Us��s��;��	�?����O��ۓw�}���J|M&�|��W�O58��h�x����=h�|n��߯�ſ��k�,����ƃ�ì~�)�������Ho҃��x�9�����?ԟg<9�>�[5zf��kś`j�C�y~��cvZ��x������k�)�ǳu����#�<���s�O��7(�"�O� ~����C���5���9=��������f�������D߻!=���������1޾�����B�c��l��˳V~�?��*?��s�Y���|r�C��;����Z�������*^<	|��:�z��꫟WH^��u�U;�W��V���F�ޟ0���Z�Gz��l�e�QK�y|���Z� a���3x������j���Js{ѣ�y|����J���s�5����������g�C�'P��gD�5Q���ǟ�n���EM^L����o���VyO�F��L�~�J�~����%*剟���>}&_)���7�_��k�ƒ��_�~O�߅�_�fy�koF}���y�o1����u�g�]�f<1�o5�#��@�e��La�����>��'���s8=�7����Qȟ���k��?/����I��O�����?�e���w\��}*�Ò'�_-}>Q���N3����~���e�w�4�11�Ǭ���ǒ�H�Z��̿V��K��s?����_k���*�n���U�_�t�gx����m��>��o˿l&��<��?�yIz�=���)��;G��y�ޓ$?��z���W��/3���U�_���O���n�|py/�t���bƟ�g�R�w������ג���J�i|��zl>?�h��}�;�������'#?�����������?����c�:���|9�/6�d�7G�?��!�����*���4>>�,��雭�~g$���p?���%����m�_�>�/�'��=b�v�o�����}�?�[��YL��Y��Rߊ��K�>����pv|���]�~3����%K\>1��n�����f��9����Y�~���Q����>�#Z���'(��}�~4�-���G��8�_-���n�x_c���ڛ }�����l�p~��׏� L�ߥ���3^u��~K�c��'m+��=�������z���>��p������6�j�uz��d�G:~�P�f?r��,�m�|{���v���g~p�_�����j��l_�h/��#��}��F���o��=�������Wk�h������T����O��_����?n��5���-r�9�ɿ���1�c�UK�Vd���}�M�o������������.�J���G����΍km����ۄ�ס>ǯ����8�N�M���yi�|%���n���������;k5�ÿ���߭�����/Wz��a%�z%�9����=���`[�����%���`ޏ؃��\����������~�#?��p~�~��YE����M��#����Ɔ��s>�B:�g{��Sci�Ó��v ����������Ku���-�����d���O+>驾�#�?2?��}��g6ڧ�d|B������y~Yۯ��>����П�����O���z��I~6��EH��w,�0�����`�u��}����&�'�Ǘ㡺�`�hۇ��xb�Z��{�X�P�g����f�B?�O���Tɯ��������_`�t�����OV_׿�q}r�[��|��Kw�^���Ǘ$���q#��l�m���ay�kD�L�;`��/z�����m���1~���z���n��У_��B�a�O�?;�\���W}�a�ʙ��(��w�޲{;�w|��!��~�m�i��+|��ܤ>��e����j�ߗ?�i��S��Ϥ���{��o�g�~²��m�����R�����?���k�S~d���Yk���'������jO��|n�C�����~ǁ��w%�盙}y����)������$K��Q��E}'�A�9�#��'������~vG��5�'~�c���q�G�8�O{ׇ ,Y�O	��>�?�~o�3/�q|ψ!�~>�3��,��<��
�h�������}>�m߯����E}�?ٗ��g��?��V�?�Ｗd����>�/[Q��`�+h���d�/$�ld�g����tǓ���㭵���K��~,~���y%����O��5����=�u_�����#^��N��o�ߗ������=]����O6�_�Ƌ����h:����A��wty�����-�D�s��Q��?�؇k���>~k1�����>�G�_N�'�m��2�O?���F���>>������ѷ�~��������z��S�G3�s^������yR����h9������x�S_�t����}<4?.6�Q����Q����S���E{��KX�����k_%?�������>�ϒ_oI�g����u�����{#�%�2�u�]-}|eϢ>������+�?�o�P��ώ�������ӳ��`��w���У�B���"�{:��>�g;�/��[��b�-}���������{
���M[�H}����ۈ���h���ʓ�������|O���ZV߹(��'E�Zw��Խ�^Ѓ��&���-�~������������e�h��j��I{+�7&������t����Hw:�����W�1|?��ӾL���O{�d�P�������^��|m����I�33�hً�OA�X���*��,~����?���&��M�Z��z�{��W�|;�3>����իP��k6\߹�P�n?��������w�_��K_��w|'�o�������74���/'����s���W���������Vc��>�5�[�Y������)��r����&?�77�g�\�U�^�t�I}j�o��\o���?zk��?�k3��@�1<���~8I߈�����E��xR���.���ת��c��۫d���e���߄�cf</���ҽ\���H�W�c=m��b�IK���#�8���FM~��Rֆ��71� ��s��O|]r�Ϩ�ܵ��L��������%����?�F=[�����;.`<$y>���~��_/��<�����i.ݔ�_�=h�����Z���㗗�ޓ�_��W�o<O���=������[��H�g��Ҩ�{ۤ~��O}ߊ�彿��,~�OyIx���V�x�>I�wF~_m�c��>���ȟ��nΏ5zr�8M���ϖ�$�?���[`ݭ���wE�7�˗g��]�~�����q���_/�5)�������x�[���;�N{Ȟ�|���Qu?�S��~�l����y�;q����������g<�pk?A��n��\F_�Q�����.�ދ��j� �_q~�ƃ����Y��Q��ӓ�%\t�%��@�/�燢�1"����W���q{������E=+�m�Յ�;d��n��0>���׌g_�/.������민o���G�?�S������C��;P>�O�r����?��ګ�},��c�������i�Z�?����u+ꣽI�[!?���< bx>:��S[�a<�w�"~~ز��>�e�p�0��|�x����O����՜_�����Է�0�_��%��g!}�I��xP^O����5��]�O��-����h��?��/&�����?����_��|�{�\?j�:������C���N���K���������{&��^d�O�M�+"��ڜ����� ���->����
z�sm1޾x��"��1�Ok�(�wz����|�������?� �|t�����mf<1�w����㩳�gY�7ϯ�t}Ls緒��M �L�֟���1��-{���U�/���0�3b8��`�O|�d����'�~�W�ʄ>j�����z�#��/��읻 k�_��.Z�=�����Oh e�<�O��J�����)��Qd�%���ַ��C��ޑ��?�{����i�vٖ?�����&�����2�����v{�=-��߭u���;jo�^�O���bx����K�����>vM��d��E<�K����߃�-��H��;�/����򓿨o���8���o��z��&���e�l�7%�Q��E�|��o_������5�5w<>��#�'Z����#y��Ο�h�87�����k��[�ܿ��`�W��R�~�8���<����-��/��{��?��*�7��+I���' �$�O �9Y~OL�}]���|�4Xg�~��y|�=)Oy���m���=�W[�@yⳀ����J�u�7�)�s�57�~Z��ޫtx-�����>�o�wW.�syA{W��������޾^���݇�J�|�%y���}1�y�Ǝ���:۟˗�(����oO����t�J}7[?��]A�*���	�k-��nI����x�������ο(/v��_���R��⅗��|�������?�����@y���ϫ��?�y9�Cu���}'�V�חEK�;d��-�-�Gz�`�_YI�k�x){�M��w�w�C���;������<��o�������}H_��|e^�j
8�V�����Z��;������dS�����K|j�6�����K����:�s}����?��M���(/z^��Q�o8,���I���/���ћ����@����0�!���E_?�����>��~d���a�G����Ї�DgG{����By��5��N���u��!��>T�_��ۚ|ڇ�~�����ٌ�������ף�^�<������L�',[��g)�g}����[b�����
?��?��C�_���/��I�@�w���%��^0Ey�^�� �T�����l�����P�'��	�W�t�r�����g��v2��߲wP?�����/�/7�U��|/q%�����[���o��W��y�Ì�6�q�>�G��S�����_,}������7��	��_�DO??8����_�g�'�gf2m��:�p1ҏ�)|x�v7�'��駷�>��GX�������$�'?��x;>5�;�>�#�[��U�_ܟ9,�M`��~ϯ�x{����}M�{L���_d�Z<
���g����j�;_��,M�;�O�j��>�zK���>SP~i���{��e~?�[�:ɛ�ׇ6�?��튡�<I������q�G</��������+�ũ����p>�z&�um���G2���Z��%�i���O�AO���c��5y6���-��`0�S���3�p;0G{L��ьf�/�,�A~�?H�}�?�֧�|��A�7�e�{-�}<[�|ߊ��]�_�K�w;��G��P��]��?[bx�2M�?�ɱ��
�����oM�џe��P��}�I��;-��~�$�����n�����=-���ҷ��{ѿ@��?\�T_�O�/;���>-���paR^��?I�{5yA�&���ῑ�8=��5������ϑ�<�� ��u���w��'?�[���s~�����-��i������G�?uv��C�Q�߳����Z�Z�/��y��+��Wiէ��#�t�/�׋�߃����{�`����m-������<χ���_�7���)���/�^��ߵ�囯?����=:�Os���[b�oS�e���1�2}T���+��!�?\���^�^�[u�5��D���{����	���ׯ�v6�	�S_|?��H�w}��}ю�[�>�ӡh�c�_��9=
o��nd��֓�z��c�_��"�i/�?�ק��=����O�x����a忞��'z������<��N{	�kv7m���������ǖ�n���?G�;|<(���#��+IZ�=��/T�����n�������ޞ��o��,�=�����I�`ͅ�>BM�g�9_5��{4�G��Ǉ�i��ҩ��C?��������;�y*�_��i���3b�w{�~��Jz��)ç6^Ģ/^z�2:חk���T����M��?���Ivx|Q�~���MI����[��p?��f��Y3y>E�?����˷���]~F�{�o:�����+��<�q|��Q��}�l������G\�	3>�d�!ͣ���Mއ*��\��6�ؤ��}+�ϡ�\6�[���1�ɯoM��O��;����{'��f{�ɟ�~Q�oNֿ�@:���J��?C��O���+~��{�'�����	�y߅�'_u�}����?�e?n���=e�����~.o�����}�4�S�'�џC?��-��4�㧹�3I��?��i���i���y�����M�^��O���t6?��T�ӓ����zK7������G�u>E|"��$�l��D­�i�.^��o����O�}G}�m�.��˗�����-��#��Z�ה����h�_���R������@����>��7�+�{���x�������K���/�h��A�@�|P�<>����0Ǉ��k���Z�~|r�½�,'� >ˀ�P��}v��������.[��,�O����c�������C�;K��O|ݾ��*;�d����?��_�~/A��3�]�ҿ:�?-z�:��ާ��s�?�y}:K��9�[����g��D~��϶��������Z���?���Y�_�wB�7�G4���/e�'����/����${�L�?'6NO���$�Y�i���>�� �\�.�?%���W���o���G��\������g%��oҏ���:��~�+���
�<������;����~_��~wS�\���ӟ���}��������������e�-��y�B�?��0�]��Az$�~g��}UA�m�W�;?S~�|�f�ZI話��D�Cn���'b�?����a�O0����0��������'ңe&ӟI�j��
=ޅ|I��Џ���??��D-�������u������U���O�}I�xOi��[+�h錏L���q�]�cs�K�s���-O�\���e�������b���^��n�;�}�����o�G�y��?�A�w���~AK��j�0�_
�3�vD��֋B��{e��~�J�*�����Y^�{S�/���~m������?l_��{#����o�֕?��j���C��x�^�y�oD�~��ڏ&��q�ge{���F_^=fV��c<&��v�8~5~� I)VϢ�/�����Ǉz�.�u���}��������睨�����{ϻ�|+~�!��B��Ƈ0���VHg��V�^���"�{�N���W���x{+�/)Yh�{�OP����5W�+��R?�{�~�Y}s~>+���3�/��R�'�Gv���D�kś?'��[�F�͉�ӕ�[����_��d�����}<Z�#�ǯF��|���+����8��L�����c��uh����	km{`�_���D:�)������������g�z���n�{�t��v>�钝�4x���:���V?����0�w��|�n�ojk����,%��~��YI/���w���j�_�����t�w,�����E:���H�}����-���7���x0���f�I��k�W��ޢ�*�[�o_�y��I���o��?�������>���ͻ"_/"���Y���;?7G�$Ϲ?��/�Q���g�]�̞���Zw%ڧ=5b}�x\��;^���S�p�^��xI�d�5�O{}_ϨГ�s8b�?�,��O��'�O�<\/��2X�����ğ������I�}�Z}|O1۟������4��sx��1]��@��F/�7��+\~��ӣ}�r��1>���~<_�����?�կ����?^ˀ}�2-��'�Ip}���߼�g�AZ�_��?�r�l��r��/��g���/���sM�.��^��_�_(����K�|iOh�?׷���������$��tC��F��o���_����<���a����L��o���h/�����_�wv���8V��7J�y�㫽c���ވ��K���w���Yc����?��1I����c����g���zh��z�'��?����B�)�2��}G�<�{yٞ�I}�����>d�j�m�72���_�?��;~��o�����Z��d0魱��9�玀3}l#�����}��d�����lN��g��6�z{w�߯b�-�O%���ב��5~\F}~�,_�1x)r�f��< =௣�ۅ?���ch�~����e�^���S6��>�o��9�����C�?km}��U�}�o.U��v�M�����o��:�h�o�ԧ�q}pZ~�2X��S��~�|��<]��z���aԗ���?��;�?�	>5���:X>oH����cOR?���5�-��l���Z��������q��/���>����KzL���܏�����s�@~٫�?U�s{0�{���p�������;P���%��Sc��<="��.e�O,��x��5}�u>���[�oO��ڎ��[���g�X<�ɰ,}��Ey���S�����ۡ>��pA�����89ZD���q�����y�N�ǚ�sX��"}��V�����ӈ������M-�����U�}�$��/����o�*n���l�^�b��zJ���L�c{�?��o4��ҷ|����oD���"��(O{J&��w��i���x �����}E�.��V�0���+Z�z�+���W��������c����Ϭ�ߧ@�l}��yl|����g#��e��_�n��/"��#���0�}-^��G~��G}��E�������ߍ��z��?@���c���[����C�/�WT���O\/O�ȃ���4~��^�^?���|�"�����qګ//�_Y�����������%����O+���kkS�`y҇��<�p��1�_O��V�]?�L���y�Dy�Xs�f�x��Gş��;׳�]X7������W�؏�-}�5�	���?�����i�`����G���ZC��?���(����e��Y������"��#	�����+k1�/�#}|��_�/m��`�ߏU_�_��N}�wR�p�����f|t���l�����L�֣y�3�~آ�����O���A���4l��#ܦh�����<~9�s~jn��vk<ū�G�e�O�8�&���<�M��G摏������q�맒��X���]�]5�di��ę��4���!�����'�/�4Xc����&�7Gn��ٿ�/��e���|=�����g���E�3�����,�x�u����g�MzR~\T��C}>~��;c������?�GDO���Vm?�������@�G����~�`���1>Z�h/��Q�w&�7�z�5{��E��O�U[/]?����?%�O����}E��ҥ��H{]�WM������Oc�߸�F�d���_/G��O�����oZ+����+�s���T��9���i�k鏷����=�}]��x}�[nO�|uy(^r���W�ϱ9���}�	�L޷�),$w������J��^�����菟�����w;���}+�����9��;�����U�w�_��M��~�n�͠�t�&��>�h��v;�{< ����c����w}�x������x^��T��5���<r{�B��>I�~�������z��.�l�܌�8ߧ���E�^��5��'��?��h#fa~��3��������������]����p�E��C����Y�_��~ߐ���D���^���vԿ��s>g�2�ҕ]^3~ޛ��oО���� =I?�G��)���W�����x������E�>���G���7(����n�e�$�|�2�~��������p~�������f��4�'�t�긽D�J�I���Zo��3Mʳ����e/����Js�����;���P����o��B���y��W8�S�~(��x5�zQ�_k��G���������$�,����c�_��o���"�8=$���j�I�xϒ��h�K�ȯI�������j��������_�/�?衹s]B�Y����s�.��_������o
�׫2�~^ �|)�g�)O������u(�����c�ӓ�w�>���>�����S�rzhn2�����9b�����fԗ��!y��Gj���k��?���[�m�%�_ӟ��"��-������#b����S�W����~߯�/���Gߟr�����%H�ل>�ﬃ^���g��3���2~��G{]�>KzE��T���9Hw��ђ�W|j�]K�g���d��[�~��i>�$�5.�ߊ�S��О�ϕ������(�3}���� о�6�cd�Y�u}���9?h��������?�e�����~���?��j�g�R,�t��zE�3�G:�3�PYz�*����������p9��;����n���������>��]�����U.���{���SP��IO����-���)��x���������#�����/Yۏp?׊'��[K�W;�d}�����/YZ�G&I�_��������(�O���s�������?��yy��Q��h/{��}��?�최��ܟzy�
�x���"�O�������z��s�gz)���1>��e��7����G���lqϡ�?Iz9�+��)��@��{�?��[�3M�ӂk�s�G���h>��O�V{�;>��˻����y�j������}n�!~⿫��HO����/��3�&_�sc��=�O��/,��I�5���s��������Q&1|���۹?n�˸�#�9=
��Մ^�Q~���?��p��-����8����k��i���Y|Jɢ���x�變��[�؛�?��a��}����8�G��[��7�
�`�u�`��1���?jp��r��{�>������E�,?��^��=��ђ��7���yz�����k���Y�
�Oz��kO/{��MI~�5���#��1�0��k�Ͻ���|>D�Y��7���=�t˷��x���~I�E}=Q^����z��w3`�k���?l��Z�A�Q�p|��-���{��a=]� �l���":�������\�_���R���g���N��/t�|�~}����� �Ϗ�y�J����?��2�/�����mk�z����4������?��猟
�'/D�ӏ�����7�7�<���F~�^������Y��e���Az6�����,�|M�;?�=�ע�{&�i,��1^���d�󞾈��o��Q�/@{�����/��|�9=��(ryqM���hO��_���?�L�{�; =����^��Y��o�����`�9��m}'����Q�P����"�:���׶��i߮�Cze��~|#�o�r�ӟ���-�}ƛg}5������Zo��9�	�?���.Y�^^����~����k�,����C¤�&��}k�����y��o�v�˧{��}џ?Z_2�h������KԏU��w�E<g}��9M�����T�{��	Ч_��4�y�����\K_��Y�m}�����'������}�����w�������W���4v�~گы����h_�~���|��7�O��1�/�O���Z+o��H����yA�>��������oUރ(��q}XA�������{�_�2����W�ߌ7����E��zHzq?���_�������|���|���C�ն�'�bx����7.A��OƧo�f|��h�ǎ��]�N�/oɏ���xP_؈����+��j������Q��c�M�O�!z~�g�S�]>�>C}�������Z��_�5��,��@����F�nk�N�����������C�k���{�������������6X���3��"�W����S^h|�5����ѿ�B�(��>�/�>�������П����-�����j�����������$��������wP�rX��<����5׿!�߲�#~�x�����^_��,��σ"�����煼��a����`�_`��9���@����듬~*���ŏ��8>�}��Z��$?�C�S�G}�`�E�g�ޗ��z�xT��ؿݍ�"����E��@~��W�=���y���Kio�}wFs_?�0�u����5?������?��1�o'yy��ODuVc|f8}��)�� ?Ǐ�Ǭ�a�[�]�,��s)��'-'���96^̯?�w�xuk��w�S�����ڋ�'Ig��Uz�q�#�����K:}�~�9����j�6�)�H/}�џ��\�X��?$>-�T�^���[��=-��m�������扯Hg������o�!�g�����鯳8oE�����z���-�f���-������+���4�����~�G��?��f-�x���._���~����\�?Yj�=>Q>���[F۾���E_��C{��gM�8��ѿ���P>'����?j�9,����G��4��Y��Ho_�5kh����F2~`~��׀���������~����럤�Y1��y:�ò�d��+1�o�����~�X�����_OC~�j����p_M�k�y�^���A��y��_D|x���}�]k�S���)�3]�m�x�5���h����R���NC�Z۲�zڻ\���>������_��+����㤧����G�~>����~=��eц���_�o~�)YD�6�O�}�ڮM����ϲ�O�^ ���@������?��&߲�S��z/�������	�į%����r�`�o>�`�7�~�>�����\�x����-ޛ��v~��?���L���z�����C�|��e૵��7�>�kȿ��"r~������O�f��{��u��5{sv_Cey����5�/��Yښ0�������0�������[�}��8��5~~�pIɞ�g�{<���m�h{9���y�S	~f���$/5xw��%5�y�u*�`����<���Gz1����h���*p�P?�g�~Ay���Y�o��g���:������.�x>В�5y��(��v����K������oF�� >3���3v���-'�	�u�����9�����2~n��~�W��y�ݢ�~��5���[��ڣ��?�{��A�	�鏙�S���Z|�ː��y�����N�<����U�Y���~7�o��}M�;�M%�ۇ9�������&>��\���z�0�?��<����w��t��/�q�L�����d���M�\D����I�W��\�wƿ-�R���W��}���~���������������k�"��BX��f�#���/��UO���;�iR�6^���y+�g}��%�k�s�FM�L���}����w^1�X���S�ۖ�A�Z�K�����ef��/�C?:�i~0���_��k�H|}~�7��P�'������S�7����Q��k���{�F~������l>Ҿ�t�Y�ѿ���2�/驽�[.�D�>����W�����t��I�ٿ_��|���\��^��<��ۂ'1�����O��5O'�h�q��kK�_ۂ�[�՗��YѶ_:��6�e{X���K�Ay�G�C��������%�Dy�_�4��㔧���&�I�Y���g��wE��<�ҧ1�������,�/����R�#@�y�Q����L���t1�wd�������c�g�����}��7����D��_D���L�����@y�/���_���KK?��]�?���}����y�z6�c�%����e���x��/����s�]���9�A��K.����K�W��6��1>ğ��F�w����x��^�/��K�������ǖѾ��Q���E_�߈�o ���"�e�]m�u��
~?m�-~.��S��]����}}<4V���~��թ��s����z��~��6����K��>��R��y����h�� �%�O��8=Ծ��hm��%�?�����KW�>҃���E��$���x���3c������9�^�{򻼯���g�5���`�w�q|E�I{*���x/��&�����������/�M�?��;|} ���P>yy�Z�_����_��sz�?�4���S0�C\�{:���>�]O�g��1�h��^_��{V�ӵ�Ӳw��t�˒n���Rk�獞N|k�{�-��� >3f�|�~��1�7d�0���o��7ϻQ�ۓl�{����� �g!?�[�����l��.�����ñ��G0ϟ3z��C	~�?���+���ezD���f��Η�k�g���&��K4򳿷����E����^��͂]����{&�]:��:-���o}_��L�
�Fu�}��忲�	`�E�^��"���w/�I�Ek�������v��+�_�#����Z���#�^���������[������Dﳸ��|$�.D~��/�?�?�1�?��ۖ<({��g,���$�^п��i�XO�y2��9��bh���8����w���Q�������5I����Iz����|��'���7���a�kɢ��~\�/@y���]���|?K|[��>��%I~���$�?`p����'I�yf�>_e���\��?���g1�q{��o }|1�g�?��G>^�߉�q~���P�m���Ϫ��������g��gs��;�K�>!)O���-}�F���������V�|��+������߬F���d_���m���ܹTq,��F/�/ϗ���\�B}���~�s8韾'P����.�Z�n4�����=�ˋ�������P[���x�<��ߵ��x3�������ҽ�0�t�ߎ�˶������h�+���w�����jp�^�<�<=���k��8��j��>(퓮�I�_y��Ix}{����3j�q{�2�U�Kb��z �_�T���^�>�`��N��O}��'5���)�2���=�6�Z��[�ş+*��Iy꣼?\�O�0���r��ӧ�w���_��J+>�û+�vX�����'o����ڻ��[஬5˿����~?\�p~l�?�v2�/��i�������;��'������}=`<����}||�(Y>n0��g�6������Ӌ�Q�E_~�}��?�|}>]���_H����E���D���R�h�N���)����5���-k}~by��{��xK��������������'�ԟ&鬏�U�_����j?�8���J�?�#L}��/�÷����υ.��������>�'�/[�D���8}j�!�Ǜ�����l=�y錇f�h��!�	���_��<������+����賒৵駒t���$]�{J��.o�R�xu�_I�˅�k���A��֧��<�A�=4���S�72�َn���ן˗�*�3}���Q���_����s�Nzd�yD?>fM�g�/x~*zd�a�?/^�~��O�y�K���gz������}B�xy����,Z�}�c����~� ?�w��<>���O�`�e��ђG�$]�4���1��޾po�_xy����#���5޾�k��������������n��e�);"���������o?�9�U&�|��>H�>>�?~�3��}������ssA�L{fK����w&ҝ^���5~�?��_���_���I{[����q~���Q>������{�mG���������~��~ӿ-�oG�}��p�>�u����ߌ?D�����g�Ô_�/��{�����Y1�Ϛ&�s�R{�|[�� �D�~�R��_-�㑻��^�*����O�}�&��}���������>�����}�����#EK?�ݯ����~km����/�<�;,٘�Oo}���-��G���� �O��C���1Xs�����S������|�<������(�Ozw(����+��ӿe=�����=h��)k��Ux�x��_�=0��d�%�k���C�﨟�W�����F���������gu��{�����y��>���_O�.�7)���������E<��?n��_����|�g}?��;D_?>P~/6�5��}��O~�� ����������w���;Q�>>�W �f���/��W'����罼��d�V_w��.�wK~��A�k�bv��6~�_���t�?Cy\���e��EߟH������I���>���ڟ����~�H�?�v���g������-���_�y{���o���U�y�'������W��=~���y<��:�g~���֚/����޾^I���$?��ܘ�>���g������Ϙ���#����-�w���$~�g���������<Ƿ&�\���l%�߲_2�����E����=�?������l]3Xm�<�O�Mm0Xs��3�W.K��_�_r��]�m��~x�� =#v!R{�r�+='��!��"ԟɷ3��ީ�&߶yz{����A���/\_������_!?��~����?��Z?����tғ�^ӧ�?t������]��'�Ͽ��x�����T��+��KZ�>�t�7,~ry���%��/{���%������m'Y<�?y|.�~y�=���� ��O�.�?K����>����˟�1<��p���؍�n8;�U��+���u��������A���^���F���Mf��}h�O������i�����ӧu~ٺ��%���6�f�%�D~���?J�>=�|���P{�����YM�ҟ�����:|3ʷ��h����џߵ�v��?'���4ѿ5�}=�ٸ��\�47�^��|�9_k��Oz}��!?f��*��U��;,����$˾��џ?��������������f��C~��0?���x�&��� g�����l?#���5���^���qzJ�����ѓ���^~�'�ߖ��ח)��o���|��O���Hw�sk=�>@}b&s���X?����=�o��gwq)rE����+IտK.�t���F/_9�j�����uo��=4��5���-|X�Q������@}�g-^�w��d������k|y(���U���mڷfk��<b�����!�������4����j��������So��|����_k�ˣ�bh�s|�����諒dS���|����@}</r{U�=�'uAi��_�~�3{��w�YW�O$�F�s>��i��77�!;������o���(n�����__�/�����t��|"�����Wݮ��߇����;�}z�*����k����\�b�W��x���1�|+����D���σ�����1�?E~�g���Կ"��M������Q��^�w�
x>���~�������^h{����Q��N���Lf���uH�|d{�Io�gu��p}�Oː������~��R�<�ę1|���ө��'�����>-y��?cy����|���}j��<��5_���d�U���~m��Z������D���(~����믵����ۺ/�����c����s?"���h�������>�^
�&�%������}�B�<�h���O���nu<������h���>|�K������~�����?}��C-}���uvD�O�z���ؤ=ֿ}{�#�w�^�������������79'Ig����X�v��\���	������~��)ׇ�W�5A}��>;Iʷ�*O�BOo���{#ϲ���ҝ~�A�������}"�/Hҥ�;I��@|H�i���w{�?���C��l<����~KX�yp��	_O�ֹIy�G{���7�E�y��~1I'}Z�y^��a}��>>:{��$?�[5z8}���_�}"���}5�?�t��>|�l����h�}�W�z?�	c��?�x_d�S˒��Z���������A/�# �S��9���}G�Ov���q{�i���F/>Щ�{Q�J���ߌt�?�����[����I������l�o�dB���;���{��[~���{�����a�����>Uf?%��F�l�����7߃��O+��W���?3mz�]4�W�kX��Hwx�i>^������r��<�����'����Sė�k���Q��礧�5������|�{��R{���߿:'��M������쏸�d�>����k�x3�7�%��Iw��+X�G����F����|���v��g���2�Z}��/�=�g�C����OMһڇx��L?f:ﷳ�9�������[M^n�#P��k�_��'>�g�-r�>-8P��J�/'�#\������*������Gc����e�=���҅~��s_�����yj�g�}9��+�oѠ7a�C��ڢ�&��w����-������(o�wEv,�d��ω���#�������Gm|[�L-~�`��O��x�{]���|?���߈�;�:��{`@��Iy���y���?<��x���`�{�^�ٿs��_>���g7G�_��W��c||j���+Y��C}�V��w�T�,��?!ϫ����C}{�g�MH����Wmџ=pv��*��������X�8���Y�����ٟ	�?��}r����Gu//���$�ώ�}PʯM1޿��>�� ������3�<�nD�Y�V<�����u�p5����S3>����A�~�ޠg�O���я�?^>#���Wj��?�?��no��q�����+�o	�����?Η�F���{����~��a����4��s��~�J��![��R���������(�j��$Io��U$� �����8+����EO�����_���]s�����xYL��w��y7�S~��(k�������􅈻����J}���xE�^k��~��-��
N�`�e�l����m�U���2�4�/�_�?�?m�~%�oF���"��D�ajp�������~�����*�;�����m�~��k�O��,F~�v���?�+�oM>���D�, �OM~9,��ߛ���y�)��wT��s�Y,{��\�)����R�����ԝ��zt>���Y=j�j{ {���ů�|���I��>�i~���E�I:�����"�ˏ����c1�Gڿ��Lo��5����i�4`�/�|}����
5��#���{-��R�A�?<?�1e[����'���̭���7��Uʧ�o)�%o'�m���c־~�Q����<�oK_��x~�u?�����g������@~���)�'�=�u>)��Q_k��Ŀf_�}�����^v����|�����6�����`�������U]OL}����*��8��K�� �;A~��tc�g��<gFS�ϯ���R?�f���~��f{L_o��qy������?�_����/���>����4�����ދtxg�������|��k�^^}��������������~&�Y?����mO�k�����|�z{��@k}i�o�M����mm}p���<�q��d��{����w�� �o�{}��5�ֽ������P�����?�3��f�������?��V���iO�~��F}�<T�r?`珰r�RW��>-��W���_�Q_�OH����o��)������^-}����������m�_�ù����\>�k���$��^,~��}��ɛ�~E���}*��Vc�?�����(1�g��-��?���l��܌�ݟCk��x���E�q�$�l��$������||��{�����n�5�=>�x�c�m{�������l=ZA}�_�����������>{$���_t����x��Ϫ��a��R���\�n�xߗ�G�D����|g�g�����;�?��/Y�"�c�'���ȟ��������,�>0+���= ��ɤ�����%�EO�g2���?��l�./֢�F�	~��5_$K<����Uh��OO��$�W����+OC��\>팾�����?އ�}���>�>�ߴ�W�~]t��2������}<Z���g3�/_}��Z��~���|��׋@//�%��H�+P?�W�+z���T����.ߺ�$�?�~����ߊ�J���Ҷ��/��?��6��ӫ6߳񸪠t	�;�k�G����O�jЃ���a�f2�����C���-3{�z��ݫ��lO��ό7M���vY|�����j�_��>��.���>[��>�7���[�J_��!=X��w'��������H���yُ�zB���A���{~�#>~_U���fs��sX��ߐ��K��W����7��=k��'ڿ��8}�[_c����#r|��8���U_���ҧ���Ofi�W�<b%���=�ۻi���s���=�>�?��g�~�G ����i�Ay����h�.n�(k{ע��&{ߘ���O��4�o����e��߻c��5}���q�nDlŃ����G�T�ͭOE|[��-}��������OD:�������2�s��Cu=�����,��ҧ���d�?�����q~d����Ozq�k�1��f�q�4���t��ꄞ5���d6?4��_z.�̾�������ͻ}J��/�?�/�������!�7$���$�|:ڛ�+����������O�i/�~L�&�k����J�<�O�=1N�����"�gi�oVGF�l>K~H�/��_c��oћ�ya
Xy]�J�pFғ��-���4ޫ�O���\�>���˴����������>�z_�������k�2~i���P�)<�py=[�g�%1�ߣ���,���я�T��џ�ߪƏL�x�~����5E�t�Q���3~��}:)���?��vz�?o���7���/��k�?���g�J}�_v^5��=��3G�-���Gy~����������f�b���x�2�+��������,��������W�_ҳf9��ԥ�]����>�lo�W��g��(Z5Xme�Q�"�K6>>i��U���U�é�����M��������<�{�,�������v?j��W�ί�?���~����g�?��b�����T��8>���|��|)�O��/�q���xp���+[��s�|K��z1��m���ޛ���(O:�;}��n�����o��G�Ӿ�7��.�����a��}i�?
�<?��҄ǻk�+�??���h�/;��4����O���s{wm���m��|;-��%��k0�y��+�U�uoOc��/7�Z�_���G�?�̟���y���o�[���(�����3>ۗl���|����?�A�|���ї��z<��|�����a��ʯ��RH���}�L�V�;Z�����G����l=n���>�l�d�5kOc���gn�k���|�y<L�=/����4=I_�w����>����2_/N�d_Ok��̿��Z��ԝ�^��Q~��-_�';od|�y��0N�<���g}���%{O���_��E#�����򻼕<��Wb�����K�+�~��ޯ��)zx�R�Os��彩��?n?R߿p&xe�כ���T���ǵ�-�/9>>�G��߈�������~ݟ,~�JR�z���������=D�'hه����Z�N��w��g����ŏ��������/��ow'����j㛭��i�{<~I~���{����zv��Ι<�x��4��$?��ɰ�����$>�їOLg{��5zg������?,���5�K���]�I������p�=_n���"���I}�ol�@���^�׷X�k���n�u_+���������8^�M�W9�=�X��籿5�?���By���<j�'�~�`����kP����I�G����V����z��ï��7X���s�����K^��X _껼���y<H����~l�����)_�ϰ�����Nі�d�@�+��E�-�y�W_���K �j�aڋ�޲�������\=���I��Gy�����k�J�'}�wz&�;}���5}��Cs��_Ɠ��1�?fe��}�c|0�O�4�>N�0�â�Ӓ�8�4ܟfg��\�?;�#�����/�g�݇�F_>0]�x�݁�qz3��~n������֟��M�5y���ü�W�;���m��R�r}��0֞�c������)���~&������9�+�i�����b�M�Ǿ��f��,������
����E+ѷ/s���8_Do�����/�����ܯ,'�
�S�j�����yAR���C�OM~�H���I/���	�����ܟ��>[�(­�������%���|r{��r��������;�u�O�>Y<�e�O�ݼ�kNb|�������_���Q��z��Z�����:\���gN���|��=��Ok�#�gw��.���[a}|���hЃ����o�ӻ%���?�鯠���.�>XÇ���������<��p��t}�B{�l���������Dw�2\_iЗ��}T_o�b���&�Gv�ݛ���>>�+����������֊��g�Jʓ��b���K���`���o���Wk﷐���\��!_'��l>������si��͚k�����L�+��q�+�EO���B{Ok=�~��O-��G�~p����|��1�-���xb�o?�`~O��g _��?�GΏ����q���?~?��%��I������i��M1��L��� [����ݩ__���i?�]�����ԷX�\����/�w�R�7����'����৳�M������3�5{0�s�dۡ��c����8;Q?�%�3}���g���#�~��G����	�/��k������~���[��޳5�������۟i�S�I��?��T��3��@�kv_@��y��s���`�?��K}E����[�?o*��G��q���P����f�W������o����<ӝ?�}/�;�7/A��׹����AO��O.@���&P>�)��J�d;���� =Z��Z��=�߯�ٓ(�9��-��Iy�K�������;�;?k����m�?oP�f��h���!5��c����;?��5���pw�����s��^k��M#��M{��_ ���{�{����?į&��|L}w�n����Z+N$�d��o�G���g�{�&|��}7���X�3{
���6 ����f�x�ϯZ�Og��Ϗ�O��������_���v���������ۿ�&V��?��?�o�M��	i�a�h퓾�P_v=�)�����J�ނ�l�\_�T����Z���$����Aƣ��R?R���"�K����x�}�?���<%���M��k=i�K�~�����y���
��A��2�O����-�|�(o�+c�p����k@O� ]�������"�����Η�F{��oQ��>�+r���_���'�?�]�ǳ��� o_{�7�>�k�=�۷4����(_H�������ї��3�+�ï|,�xµ���W�d��y���Wi.�0O��|O#P��o�Gڧi��F_��d����#��E�H{�L�q�|�q����O��%(��O�M�o�|b{믥;?Q���A��oh������UY�*�%�_�'���C�H`��=�sX����#�k����,��}J�� ��U����Y�G��7���Z���H?ϯ���×<���ꏏ߫�������%_ܿ���y��.ߖ�W��
�y��Z�N�K������ߞ�W������O���'�8�S_�.���0�ѱ�Ʃ�ͽ����W]��/*�{{�;�A��ߑ���غK�ho�~����Y{���������z�j�7�-}:��[��G������6�O{���p�-��|;��{����ϗ��C}���o-��`j��x-S��?W{���o��Y�����Ky�O/��Q?�o����O�6_��'��_��pu�gY�6?�`і�$]��I�K�{F����3������e|z��ÞC�/\]_���}�����GW��ҞM}�;Jv�om�/��Ĥ?�)j�$��O^QD���i���޷�z�y�8��y�L{��ߵ�7f2pl�j�}>��\��	���!M>,��q�Wc||&h�u?$�Z:�������ֆ7%�I?��y�&�s?��>�<a�������z���y��t�������M�#�㹽A��!�jRaɯ�G}��ȟ�b�}�·'���vE�O\��w��~N���c|����Z/]�L�Gۺ_M|#��@��cy��Z�~ڟZ�Rd|�g��|$����������o��?����������=��2� L�_G3^�#���/���ߏE<��I��yK$�#����R^e�]��_���W�������.��(3�����J�������w��Q���>"�{���#z��y�2�{�}��>X�_�g�����x<�E�٦�?J��f��_G!�����F�.F�)�S�	�������6?���C�q�޾�IZ{�ϕ�������7$[��}ڃ}>MQ�>k��-�/��Qd��/n��z/Z^e����򾿠�7b(߹�_K�E��F���Y���w�Mn����p1r�i _���G8^�bf{�5��$]��^?��w��X�h��Ms�|������#�x�����1�'�)���>~������ߌ���{��lpy=>����kmr{�_�������&~��+���W��1�`��S���&����\fk�χ,����x��������{z�o>��H����Oc��$]g>��U�D{�n�_3X�F��g{Z���}~�EVv��yn���l���"����c��U���Cy_�y�T��[��[��0]c��}5����d;����|���TV^���q��j�yN�/���/�%�G��o����z!�!�Z������}`�33^�G�<?�,^���?��s��J:���c|�y������}}A����H���Y_��K�35Xs��o[������k�E�ߒ~�e�k�	-�j���}w�e���7b/'=�?���yGm�\����>�-��3~k�D�_D??_h��\?�������	�)�j�`����?���+��/��P����Ezv���I�Z�����.%���"۶���/�&~��z����I�3^5�#b|�k鴯���;b�O�:��v�"����1ю���=���t�7k�^x_���_����O6�T��W�Ɨ�=-�1�)����z��H��顳���b}{��j�P_އ�{����k��;˻���7,�p>�ߩ�e�]���$��e����p�^����y��l�x˟F\�)K���z��l|I��Oڡ��޴C�w���3�*��G�_��[��7��������4?i������_cG��^����7�|� �����0��>?��5��ѷ�/.�4�|�\�ܞ^�/S�y�5�g}�t�wʛ�D���S'1^?Ǔ��m��OM?���7���{_a	�'�G?��M�s8��1��Smg�}D��O}���O�m����B:�M��?o$0�Ox{��!槿=�[���瑚�>^�����w~��?�t�G��ߏ$~���O�U���2>��RI�����i�=`���=Iy鿼����GK������%Y���j����t��=����	��?��b���ɋl}��7{���v�F}�n�;���5˯���:�Ϝ/�fk��Ӆ˓�O�/���_�h�_��/����wj�ӟ��C����#z��J���&����{+�ğ�5���d�U�?���My��oI_���!��/�oƛY����5����Jy�f�h�d�����A�~M_��c)�$^i�x���2�8�ك�����_�?����I���~��3���C_0xw���x��M'��-��3�b}-����}��<�yo�?<�fԯ���x�cVg�~�~����{#�����/k��_��ݨ/��,~���I��oL�>��C�w��8}%�x�{0�=ȯ���ܾ?�{������~���+�M��~h������:��jM?t�@���c��C,���)�u��=�K"�=�O����g�	��I:aҏ�l5���$���;���/�G��w������D������������'Lzi�v~�}_�������?(O��[_]����y���B⣾����������؈���Qe�xp-|����F��4��������q����������z���֋�I�\�E�S���ϓ��V�������o���>�_����Mk��o��?��YE���}�<#�������������=��>y:�������_�~z��م�󽬖>\��l�ҏ�?��3}���Qy)r}�?���o�����җ��w;��Շ5֓�Y����M��_��5;��}�$�]��X@��5���o����ϭ�ʃL���۹�?m����ˏ�Mv���|Y���E��x��/%=�_��0K�y�Wܿ��n�e���hw�$}#�(�c��'�k�d����~Rs��K�?�_�?���c|�����(���L����K��?��j�sXk�]��u֑�c"?*��C:����f�	ħ���iB_�W�V���Jϋ�?�v�1��F�_�>z���3��s�4�|���&=�8Ϟ<����I}�E�ҹ�<����zIBϚ|ٕ���g��F�����g֯����޺������Q�����ܯ)~1�s����{�lƣc�)�tG~j�d�S숾�o����>e���k���M1��1�?�����xc���s��|��4��[�c&�7ʏ��N/�үJ�G���������]T�_���忲����]_�ުo!��p�w����2L_5X{�u�3������8�� K6���{P~�xb+1���<�+��C�_g���7�>2�N��	�W:�f��|����W��ۧ"z����e�p��27:�Ӹ<�<����k�l>��d���x����Ǉ�ܥ����'J�;�S������L��}�'��G��s�>��<^X�7��%�`y��[�tڧ[�ۣ?���D_�o�������(�G�ɼ�z�~0��&�����}����i����o� ���g�5/N�u�rSB���=�����%�R^8��ߌ���w����å�ԟя��8T��	=�v?����_����$���'�[����G���N����-�����o.Y��ԇ�>�#ǫ�?@�������b}��~BgQ�We���_�Ox��_˟h
zJ>0x�R~��L�Ay��~^�}}��cʯ��O�|}��ﳪ��P>��O~�񠯷�����w���W]��Ip�[����O���X�={�Z�_fp���މ����k����̾������n��������O���'����h�:G{��"�C}��������!�������6ο�/;#�W�}�;Y���*�#Ly��Y�?�s�I�����{����Ol��|k^����]k���W_���w�8��s�W��?�6X�yu��/����o��|�Ng�ί����h��9I�,�������H���G��?�G����xF�.�$�]B_�o��<���&��bh��^U���Q����jO��q��W֚�����zh3ʋ�3{�/^��"��)?Z�_´W������gj�8�/���hO��k�1�?ڿ�:�����Ӣ}~Ԓ���Z�}4ɯ��"=����>��́�k�"�&�|")�E_���~�{����k�o����K����F�l��?�C}��![�9��~J�u��F���������?�)���-�|7����Q�yUw�3&�_������q���D�}m�޾��L����^�M�d���=��J��w�~��Oѕ�W�?/B}�-r���z���^�J�������;������7���*()_��'�&�5�w>�}"��|8������W�{�>-�l}��</��U����oH����w�sx�*�ۋ)�������[�/�Z"��������O�y���8�b���G|���xw5���$��>������A|g���׬�pya���Z�y���o����ے���K�'�Y������=]�q$����p}���~��64�=�F_�S����pw��f����+�M��D�G�'�޺�]��y1�2y�4�_����l�;�[�=n��xx�]ϳ��g����������[wGy�O���xS��������ό�����������������k��xl�$�_�a�������|�b�_��#+��������t��s��Wx���w��~�S~�� ��$]��H���?�o�j����;P~~��x��1��~��ޤ�w��l|�����n��?�˷ރ >�����x=n�[+�@yo?b��rX�]O�������R嗓�9��|Ꞌ�y��#��0�Y��=��sj�#}�}ђ�������~MoN��I����o6�e��i�����$���_���=B��}w#�������=�|~��wD?����������<�{ؙ<���e�/{/�ƿ>���w�Z�Ώ;P^���a����QI����L_���ks��_�駺2������o����J��zK�^��?y<$��fc���L{�3�4�&�Y?�?-!���t��31>��՗{'�-�Gz�~�˭	L�o��Y>~��^���Z��|��-���%��G~�w����N����f���?�|0��O���Q�L�n��R<����(Y��ۋ�e�|���?j�哭w�����{8�Ǐ�a����L��	���zy��J��l������$�a��������ρ�w����~Z�ݺ���7�>5���>Y|���~����?��F�����������_������Qn�P_]��}Ve��mj����?�4Ig��9���m��o8�y���x}�/p<j�+8}շ��OW�f˝P������c�~���鷂��?��Ki���_���t7���c|Do��ʎ���k�o��͑����V2~��+�W���:5���K��෻Bo�Ǽ�G����|��_��[������%�n2���9��S�-|��Z������Vˀ��j����j���+�轿����7��,�aΗ�}�F?ʟ,�H��ֻ��{�~V���q\���*��e�^���k�%ɿ}���^���Ҥ������?��y�Y�S�3�{^����o���c|�%{�=���?���o_�+���e�R���Fy��5?�G~�����xim�2i�������6���e�N?��7�Q�>�6#]���/��$�����:��ǯ�?l%��E�7��^�g���.[��/��o"���+Kv���]4^_�]�;Ѓ�"=k������"�&�y�H��E���W�C����^ķ忨���ɢ_����q�Iڗ$}������y�����������%���/;o��h6�}���僥�k��s}8��}�|�����@{���ė�%���}���ߏL���ɬ���C��K<�������S�d�a����t�Ӗ^d_�3�I}�����Cn����bx���_����?_l�Z��;�>����[�?Nϖek*y��9��,~��
�ՊK:o�^���y>���݇y}R��;��X�y~�ك(/�>�\�-�����ck���K-y��o����.����uK�������	�}��~�n��\؇��<��i��5�O����g��9��m�v<��=����������-}|�]m��'ߊſ��~�/�_�?�a�p�l�
=3������xuџ\���
��y~hO���/��Ϛ����5�ua��/�����I~�7���/5�����E|\���[-�������)��#������w��������w��ZO��>���o�q��_m������A~����
J���x�^�����#i�s�$�}�O���؆�ٻ���Y����z0�\��f��~sB�E�?�������jR��_?p������#]��ˊ������jA��v�~˨��e��i��@~0�{I)��A��笝d�/���|�����?k�����ty�_&�p���[y<�=\~U���1����[������u����O =�?V����o�|�Xa�Z��WV��������9}K����x�83��`�W��q����=v���v,�r{�r?�e�Gc�ޠ�_{k�G�����d;�85�?�|��O>�G������S���7���fOz�g�_C~����S�rۤ>G���+��lR~ڣ?�#��s{��u�`ъ���?�W�{��.�y��kևl�!���&���'H����^��x�-������^��o�����}֣?���󋾙�����������z�������;{��}1<���?���c����3�#�a�e���By����� ��b|<Z�7�ߣ���,Z���;�G{�������F�~r���������H���k�_��B�WY��>`p��̞���gG��Kn��#�?x��5�|����h��;����A�.�~�K�����ߙg=%����-�>�[8?��B���y�y0���	��1�Wޟ7��?�A����iH��Q^nd�姾$ۄ˓�W^����)�</���x����F<ī~��꿾�}�7���xM�펼����_��)/������g#��.?�o��|>���XD��'_�?���j��>CJ�q?����
��s>���L�o�[��G���9�����ufy��]�O���I��e�d}�W�ٯDk�������s�t�5�k�ޱ�g�5��yۙ?S���X���mP���Oڣ�MD��X�����O(���9	��k��������Um}��Q��#�׫��=5���:��^���.ۚ�����N�d;�0�s�I���G8��WV�����I{ҟ�t��{���x��2{���߯���>����q��џ�+�������C��F|\�ߟm��zrc���e�9��tvFzy�B귴/��S�ɓ�8|U����\��y��6���aͅ#K����R�Y�/)�^��Mb���ћ7�������ׇ�o/��L��4���~/����x�?��K���M�%��}�@��
�c�Ϝ��4ޯC�^�ۚ�~��&_�t//��������/`�"�����,^{���o�q�[��e����'�'H�Wn��/ў@z&~lO���#��e����נ<�Ozq���i-=��{z���'}}�����o6����oB}��5�����ʇ�?����t�d�i���Jz�|����Uݙ�?0x��^�Z녟����#���j��n�/?�����}g+ʻ�~�ײ	�_���������Iigލ���~ n�?�����{�,���"���e�d�Յ�GMP��O�wyo��o�&�?�l���'�<�`ٓ������c-iOk�Ϗ��ǯ`}����y~�c�cz~ɒ�b|�ؾt��Hg���S_�?J�xB����j�����y����>�{ƫ3�[K���/c��v��ߗ�zE���xd��o�*�1Ig$[e0���k�8��G~�}~�W�{uB�N�N���7���
���
��%h���,_�g���N�/ҏ뽾no�|p{+��^2^�"nO�I�?�ߨ?9���p}��Uu�%Ig}�'�/��@z���:���UI��h_�u��9s������o�<��u9�s�K���[��g��j��X?����ȯ����ї������G���>��]>����>E�����3��i�'����j�#vn��9�ü��������ũ���E�?�����?��M��?���o����%~.ύ�>35x&;���}y����Q�O��"���O�h���y��ˇ���䖼�.�����Gh�ٛ�^���� �#������{�����T��G���z�޲_ўX����'�C�_�tɎ��������o���e�����^�WG��o�B~�O�^��QO�o�e:�w��xj#��E�����R>�v./�?=�����,O�|��|�/��ԒGʻ��G巏o�����47����^�����KK?��!�'�C��Ӛϴ�f��+�/�{�>��֯�7��1�����{y;Q?�+����[��SH����}�m٫ٞx�P~���>��i�?�h��k�os��޿�+L�;������o�})��WW�?x}[�����7�/R���4P>���[����o��%*���DIf|o��L�>��~�����ߵw��=Ay�O���yx������I~���_��\������ПWs�훤���נ�\[�<?�g����yF���m��$��^���\���L���|�R�Dy�O��r�����Ze}~h�<
��_��k�.����WM;,��}���+z��q��_�����2�#�����	����}������]�/���	�� ��>I�n���N��!={������T�]��Z�'�O�OwH�T�����Ӌ�]����]����7���|��Qm}d�[�8�k�Io�F���Z�/���4�㵌��G�����x=�`��_��Cz�>W�o������p�$���M�~>�������W�z>�#���1�R�>�/��	�����^������o�s$����g~�o�bW5�w��վ������g�Œ�OJ�D��Z���e����ߗ��dq���g�]�o�M��g���W������Ծۇ��������g�����B��t�G'�?�y����>G�A~�������z6�z��BO����F��&?Q�c�?����q?����^h/��e�ĩ�r����Q�������t��4���gKw(_�9� �����������o_�~�4X�S��r�g�g�O&~�4����p}��?��o,��oI�D+گ�>�7���O��?��,�����&�k�7��]�Y���~Z���'��O����ѧZ�;9(�<������/���T���o�5M�m�������|�����ס�ۻ4���wK�ԧ(�3|	K>��3��3X����"��Wf|
����@}�gv>U�����i����Y������v���џ?���폾=�V?�ճ���q*f|Z_�/6��XV���>+I}����)���<���x�<�s�5{��������`5|��a����u�%�5���tޟ���x�R?��#����n����F?��7�ƿ5�g4�?��>�K���d!�;�;����O/���?�[8�kOR��/o����O��CK~�>&��Ю;��I?�5�'n�s��_ڛ�9i��?�t�C�d�D�����q<H�G�Z�?�|���5�A����}�����o_��u���o��%/���9s���e��k��������\��-5����-�H���5�Ik����f8e��?��E�����l�+�����9�w'����Wu���[�'�76�_��X�����+��ꣽ���\?4����h����uv����G��-}��;5}0�L���҃�M�����x0��^_�?���Z||[�\������tW_�Z��}}�X�By���֒÷��gJ�C�l?��֓��f�M�{��}Fǟ�#~�y=���O�7�������wV����Mڿ����<��}�G|�o�?g�p�ѓ�|9�	��y�+h�������oI:�e �m���$����2��G��R����^S���?�]f����>ko��M�W��B���AzF���_�����[`��M��㬍����Q^��}�ݦ�����������Gwپ#��B�g������Ë���p����kk�������5�|<�)\�?��1���kO��?��_�U�	\�_�I~��� >�(��O�X�/ɦy�;S���B�o�����&�ɏ�پh}�џ"�/����S���w��Q�R_V,?��*{kƳ3X���E�2~݈=����9����w�_��.I?�yL��kOK�]>�����ϖ��������d��o[�������w(��K�����\�9�T����>�'ƃ��_⧼�X���`�u1����C��>��I����$��ۖ���/��P��%��������Ϩ�iB�o�~�`�ת��s�񀯧��,Y��<���_;,}h[��7���eoU:��2~a��i��l���k��
��<���O)Ϝ���?yK���嵾|S���W�oF����g����W���ӭ�_���?��s���7D��D�?߀�9�]_�Z�������7�����Ek�w���/@y�v�`ɶI�K1�?B���(���gNO�E�<tVfl�`�5�鏤xH�D{N_͝s��j�ϙ*��Ɉ�~����f�t�5�;�Fc�3��W���5{��,]���������m"Ǘ���+�ﯬ���x�$���Vk}��/ϗy������퉖϶�ϟ8>�5�>�h��F�~��k�3ޟ�vwoM���%�G�8h�tS�Ǣ���h���7��و��7�r|I/���[��|Z��nG��E�_e���HO�Mg�D/?���v��'��>���K���o���׳��[j����?�o/�}�u���wk���{�{Ų]��"}��;)�x���g�r&��������?���Էj������yl|y�����t��_�|<桷x��I~���L\��?��_�y'���!���)��&����6����.F�CL�+ڬ���{�_����ۊ��gx���f��>���m�?�_��靾:��\��_M�� vz�:���6]��F�~��~�����3[���T�y�x������C��}��	>���w� �Gh��������11��/�p?��G5���	�g�j����KK�iR��OQ"ߺ?,�����OCyM�D�?��
7�w�^���F�R�_r�3��<�W������~N����Q^��V���X������(ߺ���ӊ�Y�$}�{����;Y����'�����i-f<��?�2���aL'~��ڼ�3b�g�a*{>��G���V����{J�N���R��4�'��U���G3{ͥ�c|�[���Ѥg+~,�k�Ɔ��,�t�$��������,�\�
W?o�<��n�P~{��qD}���L>q�j�o��kS���y| �/��xy��e���I)r=�Ob��C~����o�+W��P�.�=E�r0�S��.�^X>~�c�~�G)�(i����	�g���!���S��ƫ��|W�Kǣ?��OzӾ=-?����}$�_×����=�`���L���X@~�O?}{S�ߞ��h ���>�<���c�q���|�_�����3�%���ng%���q���S}.O)��V�=!���U{��F~�/+�g$��?����P���KJ�o5��ї���� ���������?�|����ҭ�xRe�}�`�-�@{��h���IO�/�G��&//K�٣|���~^��B����9��wE��w'�_O���_�o�|��C�c��L�xۤ����n���`������׈�~�����O.O�w�oQ[o�<�����mP>��7L�-�+m����c-���R������?������G�������޿h�wp��@�5���و��ۻ>��/䏚��$����Gy҃닏�h�$�w�.��K}��y�G���gF�Y~����q�WP�o�_E�K|k�qG���e���W_[Dy�m]?&��O���D���\���|�RgmG�)�u�w�-'���1�_�g�Y�-z�<������Gy,��¤�Z��Oo_��;��|���֢�����Rf��z\��g�ۻ�~Z�<^�i��gZ���h����o&���A�P~9>���K��t9�2�:���_���1?�9�>�o�\��v��y�鲞Mo)��}��4�&���g��D����e�i�IO��^����������}"o�v�7 _��/|����6{���F��_(��3Xgw�H��p����>��+�-��#����ԷX�������B��#�7||H���wp{9�U������5z:?�������C���^���_xW����+��ǳ�>�~)��_��A$p�~�ם�ܟq��9����i1N��𫥷��3�~���������?w��<����w&��h����C}�=.���9��W��o��[F}�y+��^���~�^X�3�L����O�[[8>\;d~O��yn�1���W������|��Gj�ړ�s���Z����v�#+ߒϒmg#+�v6_)$����~A���D:�������,^?�����^�t�M?q�ׯ��x��������(��K�D�_��x���<���%Oq~�}���ѷ���ѿ�����ל[�o,�����$�tӛ@_������3��^?��h������n)��;*���Z�J�G@���x���|3}Hms~g�Z����O���_�~�OܿF��F�w���E��}��/������>����Or<j��.�����?v�����e�W�ݟЧV��K�XM���&���d��*�����y��|����?�S�s}#~5������i���Jo=y��Ҳ�{�#��G�&r�'H���c����T����-�����xJ��6����ӓ�*r���H�����?k�Ǽ��=�ۣ~B}�� �\�E��Ey���0>�����������Y����������o�i�Ț�rz��&����!zm��+]�I{-X�1~�ۧ��������s��q�����^ғ��OM�Z��Fm=����'z|��~���2`�CY<�I竷�:�"\�g���h��z���{�{��2M�S�܎�w1��'��vZ�-������>�m�/�S1�F�kk�d{O.��2����,���������{�$�����\U��$�F�=�/��� �����Vb�^���J}�֟l>��ԟ=]{�\��?E���	-�N�&~�8)/|���/��~߇�2P������1�)/��Osয়��=�?8>�f�z�_'Hoŋ��ħ58>����ǯv���9����mM��wy�_k��iW�}�?Bg�Wާ�~���=b>{���k�V���1�?H�l�����������G�?��5��a��`|0����l������?u$0۟Wgy����]�\���Ϡ��������j�:>>����\���G�o��/����k����Ay�[�O&\$�k~����.�G���%�к��WN�i��	�{rҝW�����1	�߂�u?�������;8�oj�p:`��=>���y��3��������߽����w���ҏ>��o�gFS��L~���O{g��^+I{������~<8����?��d����iO#=k����,��Q��o�~����%~��w4�����3>pm?��F�|M���W����j����[��о���)�u)�I�H`���.E�*����U���i._���^U��z�+�G��g�i�Y�O�Em���T���۽1��I�)�l�!���o�|����=��R����O���{�y�,|F��n$=8�7�<��_��{����?��K�����1�_�ݦI����+��+�'�?��"�����e6��|Q�y�G�Ԓw���e������_��u�>�#�_���k5����'}y�]�w�]>�~|��#o����Y<��ؓ2���x��O{M��<���_1������+I�=1?o�/~_�5��{��[>k�o�|-c��}���T��^�3����Ŀ�L���k�4���_��2����������3�o\�ȯ�Ǫ�<�eܗ䧽I����5|�U�m��äo���p���-��[���|�����!��*��崙�i���}dB�����x\b���mb�>�5�.ۯH?5rzd��D��d<"��U���Gz�?���x��c�~�
���⛶���7-y�ɧ�쿲���!�㑕�������_�w�@��G���7���\�IO�'����N �~�`_�4��"��kя�?V#�75�lMX���\�RG��l}g{��П	`�O��5Kd���^�Go�ov~,�Wў�C��u���>�x���c�c��dO��d�R�W��W�}�~��� =y?��_�ɯ��)�s����b���|���_I�@__���*���~,���棗����ӕ���m���<��4��	�f��"�'�_�ߧ���oj�|ϲx�:/x����}������n�ﺾ��sIr���s�ɕ��}NHD���ּ�IHIB�#I@
h�
��*.R[5��T��QT��j��Z;����5Z��U��갭�	�y���Z���?�c<������5�\�;�\�����O_��,�s�ٿ��g����o����{Ͼ�W���~~���w��m��Ë�ƿ������7�ҕ/����)�/����|������>��=��� ����o��s���o�4_]ݟ�k����=�g�}�Y��^W|_tU�G�߿�|��2��3��%���nO�(f}��g��V}�x���X�����w��m����z4�o��M��$�������{��W��������w��;�|>����.��~����=�����H/��}����|�M{�x��~���^���������c�����������xt՟���V�����+~!�ݟ����y�?&��.�z�x[}��?��}�����e�>�?�������y�{���g����Y��}���C����뿶������x�'�?���
���|S޿;�����_��n���p������n�����^����ǻ�f�Y����i��ٗW=����z�||s��h~��ﺞ��f~��߾u������2�{���ύC8���v������7�7���r�A8~����s�!�[|^}t���0����n���_����x��~��D�'��z�Y�����=�%c�}������3�>������~��w����=��>�Iy�����w��3�w�kz��������k�{���|?�����?������>���X߫�������������s�:����W��~�������d?Q|�0�w��S���v?����u<������������+=�X�X����\�?Y��?F[��|N�������O?���W}�}<>��L��b��C���ϵܫ��Wߔ7�������1~�~��1��'��������x��>�_"/������]=���;�~B�����ǅ���������?�}~{��1�'�W~.ƛ�η��y�9�G�����Qߟ������������������c��S�r����#~��2�ߏ��?>����[|_�;��{7�/�lO�,���:�~����c�z��������w�kޟ�����]��X^<���|�����zf���r߷=��G�������]��>�׼7�S�lO������ό�g<_܏>?��P޺������xį�����,�/}���}]����q���~̹ ��>w��x�/������~}�?�ʋ��sl��Byk��x����~�N�)�����xq�����C9���s�W#��g����Ow�f_Z�����{����t��xF�//�~>�[���mO�w��_by��w������fn��������/��}����y����Y�����y]���gWϗw�����P^�|�������w]o~Y���oO��U��9�#^�|W��|�q��{]�:�����5^�׏��_{��w�7�!sm��-ǟ۞��|��p�^�z}~�N_!�7�j}��}��������˷���c����b��/���w��|�5�����^����#�O���>�}q��G�;뻮o����h����7����l&��Cyk��{��ϫ����Y�?���~l�؟�����[���k��b\�����?g����x��o��i��z���g}^{t�ݿ�c������k����E���_�mOǗ�m����~q}<����Pޟ��|�3~�cn�7ז+���j>~ă�ߟ������3�cԳ�χ�3�wu|O����<��o��?�=�?w��m�����.�n|��p��x�U{��W<ߣ�6q���F������G�}�>��w�W������ߟ��f9��i�ϱa�_b��?�iy���]�G��}��I�W�~��P���Ϸ���/
����~x�~�|;ߍ��n����t�y��~��~��z~`|e]��x�ǟ�~�����싑\���1����;?�����~ݵ=�/�z��=b}�~H<_����o�O�α�o>��=����s�˭�s�<������w��/�k��Y>���W�g9��p������|�޿�nO����~ۃ����X���4�C?���;�]�����g������U�e�����wu�8����x��s~���Z��P���m�}}���7���M���_����I�mO�=7�_|��o���8�=��L_^������)/�7��g�}�_���-��Q<��~p{�o�׏"���8�E�.�[8^磗������/�����y�����������g���xw|�>u�<�o���o��>?{?�o<C<n]/��oۏ��s��f��I�}}��k}�4��W��y�u}��_�G�������[�7�������q}�g�c>���~���}�#�w�����1����پ�?��+�>s���o}>��k��:Y�u?�������ߺ�,��~�����۷���x}�=~��|~9���;n�7}��|��>/滶�[�<�w����\����W����������q��]�z]>1���A{��:�\������G}��_�?��Wno��y��}��g��:>_�G���O4��ss}��q�_�׿d������^��v�>y4>�ܞ�ID��G�I��>ʋ���o��e����E��G��a����W�v���7���2�=�w�^＾;���mOy�����o]��<���_�{�~����Z����7޿��g�x��絭�������<���<m�����O���h=?��?���#��ر�x<��U_�j<{���B}>��xj��PN�ןϵ����oq?��������lߏ�_��7�����߰�����aǃ8?Ͽ�t���6�#�����|1����;��x��yy��{[������U{��c���a��w��c_�h�����Y���������q��m���ݭ�cyq>�Z�߰��|��~��TO0��<�~�h?�>�o������W=-�������>����>���������3��G����b{���~��|�[��̏������|�߶�����������6��Z˛uY�oƿ��������g{�귶_�?�_��~�����~�|ֻ�<�<����m�}>���ӛ����G��.���~[�o|Z�7������jG��g�x{�em�����x�������ϱq}_�����{�߯<u����~���B����#}�Q�w�h�<��q�z�]�7�e}��g_����a�7+?�����S�x�q���ǵ��]�.�/���$���x��kۇ��1V���o>�m��臨��s���?�w��쑿���Ǐ����K1�wǓE��x��ެ����y����z3���]�_�����=����<�g���O���T���l��o=Ǘ��>k<��^���r�Ǭ�����B�߭������x�]�7�w���y��+����z#�~�y����y��[7�ߏ�ߏ�v���烫��M���oU���������k�x<����g�~|8��N\���ϣ�0�����x��w� ��\����?�������_�ݿ�����������w��|v�����:�����%�?D=��>�箷�?�^�?7�k>�[��k"}7���"����?���ǿ���<���Q\/�����}�;���m��Z��3���_�8������x�z���=�W���������#����O
��������ʿ����~��q}���������������8>����ǟ���~��>��������_lO�����.����a�<�?\�����m��k�}~�����=z޸���wݴ����u�x}Mo�b�����-ϱ�ۗ������7���������������W���o�dS?j}�<�.��_��Ý����]��'��ob�����U{~v9����_x�G�����������Ɵ5>����c�{��'s��0��?޶�_�U}������0������������"��?�z��>�I�)彻�������ϣ�����xc�3�����}��f�����#�I������ê���4��F��ʿ{~�қ���ߚ��8����w�{��1��o��罿�����|��}7׳m�K[�x=b�y������h<�;���6ߧ����]�*�~ٌ��}�g�o�����Z�������Y�_Q��J�.�z������7�|�r����;���~m�g?p���JO�n���p���>�=�_�����W�s-o�(߶��٬o�c��`��Q�}�=��Y���˻��l<�=�y�Z�n?tԳ����e�x�i9���>�~qȣ������i|hیg���5�f{�|�S�����l������1��#����t5�ݵ�o��K�6�G<z^�;�B��������gt��ʿ�����3�ޏ���ǯǄ������~���|����}�ӏ�zW<����x���'����ߗ������]{\���G��X��������wF�]��z�~�*�������M�?�����|�������~��G=�G�S��G�鞣�7�M����~�>��cn��/�����|7�Χ���˼�q|����/_�'��mO��Z޼�ߵG��/�����;^�׎���n����Z����Ǭ��]���(������.��7��?ws�ȇ��o��xpO_�������/�X��|�������m�z��qI�n��z���� �~�<��_�������������c���q���_����X�s�OM�ݡ����m���?����5����>���/�ۃ�O�y��x�<�z�b}"�����i�？�zf����0�/���]~���g>����ܛ����>��Q�0>��������_����W��oO����_>��P�����g������k�U�'��پ������_����T/��x򈇊����/��9VD~a�)/��9����xS�򮾏ֿ����͘?�����@��8����w�y��/x�۵�����f{��ww��G�u[�����������z��x��������Oo޿u���zY?�k�������|�?�����}�~�1��X�y�ݿb9�٣������;�a���Q?:�w�/q|��_㳯ƿ?|��g.�?�g����?z��导N\�<�	���������������8�W�z��~�x2�?>��}<��<��޵�\O�����o���<�O����G7����m����kۇ�����׺����oٞ�ߙ�~7��m����]O����Ss�Zǟ8~�������^����b|���m��~g��7��0�'~�r<竕��/���އEe�o���a�s|����Y�����1k|f��`{��?���s-�g���=����oO���^��}�~?��u����-7����)��W��b�|��������r|��h�������i{�v�st��������|����c�7|��~߷���c�w�����q{{}b��ؾq��߭7�{q�8���mq���P����j��O�G��{���z����/�����[��w�?k>������y����~�}f<q����۽?\����_��~�Z��37�����ylߨW�n���~��>w���\�|}���������ls}w7?������$~~u��眿���x��u�t5>>����:^Ǐٗ��Fl�y��S^�~��s������Q���_?�����Eh��nOy�9���X�8^�k�����x�x}��w�w|�W��Ol��p���^���o���ɫ�c{��yͯ��ޞ�����o��<^O�_��?��3�o��K_>���׼7��}��x���;�et��}��l��i��g[��6���W�u��;=��7�G��w���~���Y��S���[��׆�G�6�/��G�ޮ����<x�-�o�a�+7����t�<��z}1�?�0���zi�5�g��~��S������\���k{ͱx�g�����>>������zx~7��Z��/;~>���o>�뷫�}��s֋�}�w�|>}e��m���U���k���?��ܔ������?;|?�����z��,�e�����>�|߿]��s\?���wlO�\��������[���A����o����3���|�,Ǒ7��E�vm���������\�?�:�'���|�.ǳ���P���x�s����[����-����s.���}�>�D����<�{�	����ٶ�{������O$����9�o�����hж�;��n�o�[�<���~����u<z������{���W���|?���~b�ݫ�x�u}�s?�k�_3~�o��ϣ�"ޯ���o8��6����b������w�����k]�ξ����7Ǘ�zs=��t<���?�O��e������w~����c���x?��x}��:�=Z���̶M��;�������z�d��g�����#������_�/c���Wx���G~f>�����>��y���cl�����+O�kα�{��9V�Ϸ���n���,/毌������xz���x�������������.�'ߔ7��o>�ǳ���E�k�O�m���Ҏ����6����z���oq����W���x�����?�/�[D���ӛ����|/�'�'"o}�����/����k��7\�w=��j�a{����l������;�o��ζ\��_t�k�"?�K���ϣ��o~������������?������^~���yd��]����}�|�?ws�����o��<�����b���}����|����-w�Wb�ν��M�~����������z ������;|=\��x��u9��v�|��#����a����6�%>�/���x���z�Ta���7�_[��Ǉ��Ϸ�^W��n8�ƛ�֏_~7������О���k9�����Kcm�����n�K�}���Ɵy����������������{��cݟ�<j��w��1��ŷ���[�~y(�J���z�n�B<������z ��X��no��ؿ��?������?����?��}������'/���?�q���q����=�"���Y�����|��ޜc�O�i�G�i>��?��9�����x�_��K�����V���5��G�[��;7�?�?ǿ�h9��⧄������k<4��mO�-�����i���_㛱�����������?���+Cy�����������:�����������a��.ǟ��y����ϷQ_>������/�<C�7���P�|^Y�w���u~���ӿ���雟_��X��o{�`��ף�ڞ�O�>�~�G6��&�������>�翲=�9?_��W���p<ǖ�S�|����g]���|��7�����?���W���ǿ��<j�-�{�>���#W�����__uS~l�?���h~��pǯ��'�����|���c�w�縟n���G��Q���3Ɵ�M^������p��7�����ǃ��	��[�ϱ%ƻ�����Q�|�&�����;}�-�~������W�����_ʏ�;�篿����N�n^�:_����U��|^w���w�^��;����^ϧ�����о1�M�s��S���ޏ��A����v���-�?��Y�_�����}~�������3�'��9֮�>�ֺ>��ݽ����g�Z��D��8����>�_��>_��9�����G�,�e��3��P�v��-��j|Z��;c]��X��]���ǫ��������7�}�>l}c�>�_n�\�+�_����7ߟw��׆�?�_��}Y8_l���/��~?c{��9����\���L_�s��9~��[w�������s�����0�by���;������}��u���M�c�<�_���W�b�����x��P��_�tS���^o�u[盻���v��"^ߣ����S�����������8�_�ۏ_�c�~�{�{��X�����x�����������Z��r<��{��w��/������j{�<���>)��v��>��~��ɿ��=������7ߏǑ����M�����_��F��8����X��ޝ���9��U���x�r?>��c�p�g2��߲����빚��"�?������]��_������q\O������{�yh�ǨR���5��X��|w����k�u�|�����?��[����f|�}fߏ���b{��������9�.�o��7�.��kg����_���S���%��7��~����c�߽�߯���������q�y���sߗ�ǳ���x�?+/z�>gm�8���(�������#�x7����kn>������7�)_���n<�����n��Z_���������]<;��?������Ǘ8�^����k�������\��8���y������9v��~���ܻ�W���x��_s�]߿}��4�7���_.��}��۞ޟ���Il�8~,����z�>������^�}��`{����}�]\�z�GϿs��������=�7�߯���-��U>���߯�G����c�s������9���*?m��U7��j���7�;y�����W���C}����k�v����}�n�_[�?�u|���Q7��.�?�U_�_�w�e0�>>���kw����N_��=y��}���_�����c��u������vϫ��p}�?=��c�����9��7�{��{u�r9����ߗܽ?���w����|����l�;~%�?��_��h}3�^�϶^�ԯ�K������������6/���y�#ϲ����w7�7��?}s���������7��k�G��O=�}��7��7�G}�9������#=�u|���ǬߟϞ������nO��/����|9熟���g\�/����_�����������wE�z����Om���]�G���~Ƿx}��;=����~W��������s�߻�%>���`����������������m����Y�-�ϣ�!�x�����/|>�{yS�x����z%�W�z>Y�o~���ϯ������sy^�����}W�F�d=~�_"��l����T�ʟ���W�3�ye��b�{}���x��py~z����������:|=_�޹���[��U����i�x<��6|������X�X�_0���P����=��G7��u<����y΍��r<���������p��~t=���?�����i^�����X�?}g]���y���'ί��U>�?��������b~�X��`����������W�^_�o����x�=�"<?������p�����6����{�����Uw���{^�g__כ�-��������+�k�-��i���՛��d\�߶���m�}g{6\��~��c�s���y������� ��m������}��x<���s���#��5?�d�����~��>j�|�����������|�M�q��k�}{��������}�c}�ֳ�lo?��z��������^n�_�������;����W����|��aZ��c{���q<��}�������w���Xy���5߷�����ۯo��c�}����0~�;6�ol��~l�o|��߽{�1�_�W���m�/��_>���������������u�.߷Ϲ�;o�����������/~p��v�>����\�?�_���O��~������=_<z����������,�~�����4�����}s�7��ͼ�u~����ѫ������x��7��/�?��r<���p��G�S�	��b����$���?��uW~�O��#��u?��;�{��Q>�w���?������Ⱥ?$��c{M_������_=/����n�Z�?}y���	ߟk�&|����ģ��ε��������n�[]=/m���?�Z������������"�׵=^��ph���ߏG��"?����_�/��'#���������о�c������S��w�W׷������������j{����?%϶����o~?��7�3����o����?z�x�?�*����w���ȃ�����z+ꁾ�=����w�~w��?������;��K��k�5/b��NO���h=:������z��|���~O�m]�̹u?�Ͷ���x��5^�������/��|��W����t�S�>L�q������/�7������x���q>��a����:��������w�_���ϝlο�������p/ƽ���x�|����K��q}�z�X?_��6ǋ�����ئ��]~�|g�G]���l��,���=���x��ȳo��S�������������v��z��r\��:�/���v�旫�%����ƛ��������?�'�E�z^{���x�����?�_����_�=�?��w�X�؞sm�7,��Y�������w�?�������|�h������<ꏱ���~�^��~>��~�m��3��w�^�~��G�7��7���}0�����������VW�A<�{?���z,�u}��o�[�ա�u~������~~?�߽��/�������g�<>��q>��ͷ.��m��w������������ӵ����˻z���r\�WV�����<�\ۮ�-^�����j������k�����}�'����X�z?f[����_�w����&�k����ob}c��Y��f�zc����GxԞ�]����1^�������)����Y��?�=�ӛ�{�?����~��_��3����w���Z���o�Ϗߞ������yp?_�Y�"y���w���r�r{o���/}z��N����p�ވ�ո�����W��n��]��U�p~7��X����1����$柼�O�硻�����<_�/�����:���2�����緧���9���N�+�ۘ��ʓϵÝ���3}y��֫q>�׷~?�ض{��0�7���8�/��O�{~�ئ>h�ǻ�߯����+���퇘����G�?����}n{���nc߶Mk�?��?_���u���wgl�'ݔ7벮���V�I�ߞ�O�|w��+��{^������H�.�5��n��WC�������^�cϷ/ǯƿ�l9��������3����~~ŧ�=�|f�ߏ�;^��?���ȇM��ߋ������\���c�z�k�y���?�W���/�]�/�y7|���+>��߮��l�����}귎��P�x�~�9��8>�����x6��?�_�'��w���M~{���ҫ��|aw�Ƽ��������ܞ>�������k��b�ܕ�����謁�/:�k�f�"��_�X�7Ǉ��{�����FY?������/ٞ�/���_���O�@�>w���׳��i�of��oߏϷq���}�:��v��1^_�����{���O�O�����h���My�?����o��H���;�������>�˛c�Oz�/s�����G�ӳ~��9�ίyz��n�u�w���_f�~�r<����]ǫ����x�qY���x��ߺ������_��s������_�_��o������4����b���~Sߙk�[o>����W��������?�n|�㭿���i>�Xެ�:F���c懽�	�7�w>�����^��P޺^�����￻Ϻ�=�=�O8����x�U��s����ǋ;��*��7k}�ܺ�'�ޞ�w����?��p߿����n��k�_��z��.�k��w���y��e����rw��������]�k{�x��������G��w�Q��^��g�����w�!���]��?�ss������|��g|�4��ʇm۽�|�=]O~:|>��.�Jh�z<�;B{��?��q������������r9���?���_�����~4�>�ϝ���lO���X���=������S�*�ϊ�����+>y�O��?��r<���e�ﷄ�Y���7��W�'��#}��^��h�����w��ӡ�����z�q��|s����5�G�?\�w��?ο^Ϝ��M{^�����v�/QO(��?�����������yqq?^.��^�����-�?~�_�=ڟ�?�{�;�?�ϫ��.��z�}}<��G��c}bY?��{���_̗�h<X?{������ֿS�ꏅ����ǟ���~����{0�O��������?Z�\�o������=�I��w����q|�B}���߯���W���7��.~�^����>���Ys,����ϻ��X~�O���?��:��ds~`9�����.�����r��>��~m,o�%�r�c�{��x�s���b��eG}����f�l}�x�S��?���,��n>����|��\��Ͽe���$W��b����]?���Y�w�3��߳|�5��q����z"��~���ϻ�?��X��L�ꏇ�ܭo�E��ƛX�9V���/ޞ>����q��_��uڷ�k��y���\�����f>���%sl��P��}��?1~�~>�m����7���{��?\�������D�1��[M�Y���>�,\�o?����;����nާ�����R�U�������k=��bq?����W7��'�׋����W�w�c��O_��w�7��_�d9~��2��K�����w�/��=��ؾ��zt=���u���[������+>2ޟ��/�w�~���_WzC��j�_���̋�������������q�??����k��.���d�[���ȻFd��αm}�����]�ˬ˷�\�;��[8~���ʺ;�5�8���c��]ߧ]���x����Ƨ�~����G��_�y �����x����Opu��#��Sk��̛������m�q�g��>�W��Wz�K�～�������髟�i�X����}���|,�����}���z��X�����=�����M����~*|}�1�ںޞ��TߏlO�wb����9���x�%���_=N�/޴��x���8~E����x�q{\ܽO��{4������t>�}�Nv���?��潍��߹)�u�O�|0�70��������}�v�<�k���g�|>��"���|?��ǿ����������~s=[h�����>�����w7������l����+����n�}�p�%���x�����[�����s�%���y����G��?�=���.��7y}^���~jj����绀��b���G|>��+������dc}��O��^no��Ͻ�9v����_��������~S~l�Y�8�����_&����]���c���ݻ�������x�GϋW|H����"?���?��|��=��{��^����<����m>�ޝ������������������w�yn��u��d������:�%����o�ڼ?�y��}]l��׶���w��wBy�ƃ�7?���p�}�>���e����;�����-�q>��U��g���Z�+��ٞ��������x6�ͬ��o_Y�������9�c���s������|�}���j�1���y\���ĺ���&����j�ɣx�����*�|Ա?}6\_|����/���������w>+������ �?�_~����Q����e�<����<����w�sW�Ӿ�������О�ﺟ}�W=�X�τ����~m��<�����;�x���������	����髛����=��yu��;c�|���������^�������q���������~�o̯����/��ϑO��m��[����}|j�k����l��������������=�g������|2���x�پQ���|��?������~�n>��g���g�~�����r~7����mO�c��߿��~^���|�(~�vվ�}��������x������ʻ[^}��w�>�7���P�8_��P����Q>��N?#^��|_�*���|������w[�㜿~N�|~���W���96����}4�<:���l��y�|y�>u�sn�����W�C��p�G�����翸�6�ߝ����ʏ�\��Ono��q�Cl����vs<�[�㸿9�q�vl��_���kϫ����������5?A�O�~�'�z���i\o�|��|�}��??9����;���R��c}^_������z/o�w��-|��������Ï�����,��_W^#���5�7��O���U���;}�G��?��k���P^�KN{=w��������g�������ʱ?ϱ��.��Y�7,�q?��M��C潊����P�8�̶\��Y�u��|���~��<�߻���_|��P���O������c�ߏϛ�y�S�}"��������������e������|�M��?\���
�}W(/�_��G珼f�%���G��0�1��_��O_�;o�?�{������$�~�q���I���uS���/��O�c�W�el�u�ߗm���/���Ú����|S���|�m��~>�~�r<����:^ζzο��|vx?�o=����6���P^�o/����l��[��o��޸������~?뿮��w�գ����x�~��Ɵ�Ϻ��0���-?��n8ޖ�G��}xm���w�M����Sw�K|ދ���?ǒ;����qw��#�������������Ƴ���z��h=�׏Q�����^��~���Y�w�|��8_�U�|��3�]|_������j=���p�O?�3��:^�i�+�|9�e�|��/��z�������>s����/Cy��4�����k����)^Ol�����j�-��Mk�e���؞�����#�*�.����ȿl�}{|ǃ����j�y����^��W^������Q<��{���������[�_2������z������=�s�����<���������'[���w���,�ߎ�}������n���_��~�~�j>���Ol�ϻ�͹�w�ϟ_z�|~u}�}���9W|���gۭ���o�{�5��b�����W�#����}|~\���o#��h��h}�m����p|��<������������qQ�'�)Ƴ�7�����?��Ayw��x�;^ϸ�w�o{����8��k��Q���]�[ԿX�k��\����qݞ�Gc<~������ӥ�}�[G��z��?�Ƕ��Ì���m3��~�����~��x7����Ϩ��/�Ͼ���t���p|�������у�_�~k�����,��z��7������Y��w���l��5?�o�7�k<��Z����/
�����}5�|�A�ݭo�|��7�������}M�����'�����;���p=?f{{�_��:^�������|�x����c�?;�~m��z~�����?�=�����1^����φ�|i�����#�c�������������������y=���|k}�Z{]�ξ����c|*��^˟|���g�[�#���|�xd����/��������_�=?=Go/�?zt�c�>����<w�~4��C>���~�G��U�޽��U\����~����|+���xwW������Ϲ�o��[̹��}�~�?�w񝯺�����/ǿ���?z?��������}'�7���a�]�3���}�m�q��}����=�>\��j��1����c����_��]{?ҟ��O�<���w|�Ϸ��|���?o|��x�x<c	���Z}pS^|������ߟ��>���������l�O9c7?���W�7^��y_�b{z��x��|	W�y�����nO����O>(���\<��w��f<.��c���a�u1��tS���_k���Of�}oy��C}b��G:���!|�#��8����7����L���p��X~�����;�0�Ϸ����q����|��_������'~>��?��b����7�_�︾����_��!�����7�*��j�|�|y7��������2����8���y>^�3�����.��m��j�����)�~�����.�ۣ���<���ݽ_ݶ��?��W~�F�����~���7�?}7�|���i��x���珞?_>��u?�����������m���B�q���'|��p�?>���߯�Ǯ���g/7�g<'��<W������z>؞�mG���s�u~sՋ��4�>�w޹��Ƿ�����r<�������1}o�q��|_�����~��*/��{�^�k��m�aǷٟ����G�k�uYy�ٖq=rw��p�Y�?������m||4�;�sn>���b{܍'�>~��n�{4_^��5�'�o>G~��}�O������_�m_����>���G^�+.�#�W�����g������g�϶ݏO�_|��\����O����翻�l�z���q��Uy������{�{�o�Z�{nʟ�w�x�ds=��/���BW���~�s���[\��]������x=�֧��c<?���Ɵ�����yo�{/���c����^�X�8��}�u}߹)��<�?�������W׷�7����������s-�H�m��Q�<��~��4����M����\"��o��>�w���ؕ��0뵘/�������x��_���~����������<t�g|��y7\��w�ߘ��Q{�s�ֿ��=��;��+=�u|����~�x���ω_��q�{7>��p�O�x���|�����1$�7����ū���?�����x�-\���o�{�^_��痊ߟ��.�U߻�2~��Ο����������̼�u}��͞�}ǧ���绹�����/������率������Q��}��co�?�Ϗ��������������o��/��{�8^��z>���oO��7��������>|�?:�һY�w����"���7�����/"���?ǿ��"��a���}�?�=���~�g��������\�oyN���������?�7�����\�?Q_'�7�[���>�3��|�Q��N��Q{L��I7�_��������	�������_?�~�����X/��z������7~C���d�=��d���\��0�П����Q�?}{������}�w����q�棜�/��c�Q�U�ݭ�c{����>�\�G1����|?旍������� ݿ�s�l�j����Uy��|����F��<R��������h�xt�;�w�ޚ��/]�G_M�~�����O=�^�ow���;_<ҋ{�>2�'�j���=*o=���1�G��y����#>��߱?�ϳlOǇ���s�O�����?�0�E��s���W���?e������� c���5������ŏ��)�G�����~���W����~��/Ƴ����Z���\����GB����?�ף�1�3�����諾��u�����y⓿"�>������^�����_s<[y��w�_'��-�󳟹���ǹ�#��{���]\O����#?�4�ß?�3�?��5��������5��x'|�a��~~(���C���#�>�G����Ӟ/���ۧB{\�w�=�?�K���������H�:��#e�}���������On�g�����w��W�7�i9�������}�񷎟�����_޶�����e-��v�O�h~��϶�~����y����˧0?[�������?z����o۞�;��f��5��kV>z�?�/Cyk����w���͡�#_��z������ʋ�F|?u������ϟ�<�����9������������=�'޿Gz1㧱�y��o�u�S=����t<��y��x�?�t�}���\8_�gb>���w��xA��������%����GϷ�����]�绪u���냛��x����e?���4�g�����w�^_���'�*~s8_������z^������~�qG�{�|�s�������O-����[��U������X~��	�_=�}z{����Z�ݍ��ޜ�����w���q|����OW��~�.�m�\���>��O�ǳ�W�h�-\��6��}�G���Z�\ϭ����/�E��w����7^Ϻ�y�O���6�����򏵼ȿn���_�z��x�ȿ����x�^6��(�/�������*>����=���&~~�o�~���#�Ŷ��?c����>/���wQ���<߯�Ϲ���Ϯ�zґ��?b��������X�g,������s�q|���W�;�x����j����������o��;��5�-��w�D�>�ÿ�����~��+~�_��'�#��0~�w�ܟ�=?�'�O������������/�E�
�{8�Ḅ�3��#���[8����R8����9|?���P��SBy%�_	�_B��p�����j���k�>-\_�k��Z���s�����3���;C�g(����P^��p=�uy_����=J4�h8�!�e�g�S4�`8�O��*_0�2ʈU���|��~Ī�x�M�=rl��7b=r�G��_b=J��/��k��b5Zc5^m�5��,-V�ų�X�O��i[l���b=�X�3��g����ѣ��QG����)J4�h8�!�#�ܱ�z��+��FC�����^yD�;��)�$�ؑb���c��x��sG��F'<�%ִ�B���ŎO�ም����8cg���~�{{Ƴ��,=�%:P��?ž�^�h��-�h5M��صS��)�@�eľ�b�N)����z�}=ž�R��صS�pR��)v�g�{r��I��I��I���b�O��O'��g��%��#EIq�Hq�Hg,#v���O:?�},�9�9N9�K����7��9�9�G�sC�ސ�7�@�q��q=����)�%:P��(G�9^K�=r�g��I�>���nv�}=Ǿ�c_�qq�c��q��qq�c_ϱ��87�87�87�87����B{,4�G���'�;�sC�����_b�/�٣��F���K��%N%��W9%�%�2b�.q�/�'��%>Y���)qn(�'����G�G�{r�=�Ğ\�sC�]�ā�ā���qK��%���{r�=��q�^�^�¨�a�ƞ\c?�����Okqkqk�5v��Z4ċ��c��xk�5v��e�K��i����5L�cr-�q�^�]�]k,4���z�}��5L���5��x�k��05�5���05.Yj��5��{r��t�]���F�}����-.7Z��-v�;�Cp�������E�cr����-:P�Ԣ{��->����ڢ��-�-���z���n�b�l=^K�-.Z�tg`�8��q%}���Wg�g�g\]�quqƮ}Ʈ}�G�3��s�g�=����3.��ؓ�ؓ�8П�'�qY|�~z�~zƁ���{���3��g|�<� }�A����k�3.7θ�8�r�}��k�3�g\�q�qF�8�Z���aθ�>��/f��Qg�{����G�q��сz|uӣ���G�q�ӣ��.���z������3=:P��ң��8���R�сzt���G�ݣ��y��az�W(=zC�K��=�G�SA�������j���������q�ҿ0{|���/�o,~�����R���;_�B������7���_Q��ue���9S�Bk��Pr��Jɍ_}����+���JO�|r��6<)�s/:�ꜫs����>�����&���[c�c}��S�`9�=�M�􍅳�{w��8W�J��{��xw�̹2%g�+[��Pg��N���S(�R�ʹ*窜�r�Fɍ������~r/�����s��}�S�Εv�7������s������s�����p.F��;����o�o,�[��|�H�<�bN9�7��7�؟|�`�8�/�⹨�s�;o��o,�!�s07�	ž��uf�:NZ����O���f��;z�ab����sS�wsS��v΅%��M��|'1%|'��$�)�;��*��J�����_$� ��9%�	�H�ś��mȼ���8{���Wޔ𔄧���~��L��w�L�S�w2�Nƛ23Q�w2���_d�"��u]�/2sJ�S2O%���2��M@����Y�e�)���<��̹���/3eV���ޛ ���+3^��ʌ�ef�7��/X���l��ef��2�_��_��2�����07概Vq�*�2e�>�WaN)�)�)<f��
��_�*�M�+��
W����Mo*�z��_ṩ�MO)xJ�S���`�w
�Wa�*�_�*�Na�*��
�UxSQx"+�^Y�������U��*W��*sS�)�g�z���x\eF��h��x\�S*~Q��*�*��*�R��U\��Wzo��V�j��Vzfe��<�TVV��Y釕�S�?�USc�o����q������ ����{sA�?7������j���Ecvh����轍Q���j��Fn��q���k�F�o���z�/cx㩤�)�5RcE�𔆧4F�����8���8���3~ce����;��;�g��:񯓧����M$���s�'3ȉ����|q2_����Z���N�Q'��ɛ���o:�/N�H'+�O9񔓕��|q�'k�/8�'����I>��<;��2�>��󝧉�t�|�?wf�N����N_�m:}�3�tf�N��� ����;=���;sJgN�� ��3_t�w�:��Y��;���;��c���Wǿ:뱎�uf��,���,әe:sJ�+;O
�Y�����܎�v����A�� �>,	K�rFK|����_Q���B��sʰd,�=��T,�*�놅+���a��8�g�����PN\�5�7,�X|#=,\E\WW��B}"i0,����{p@W}gX�O|?v�;�Wp�P������Ύ�����cǎ�@#�4±�y��㻸>���[�aX('�qǎA{��g�3�Ep���U���"8��O��lu��)����t@u�/�x�c�/�<<�q�u�A��8�����\�%���a��J�� ��p���B�q�w�2}��#������w��`N9����b����p������b�8��/8��8��G\}G\YD폃���/��K<�������b�G�O�G�S���������+�M��X¿�����&x�#�M	�I��R|nZ߁"�'>[�Κ���+8�
(�a�d�	B��8��Œ�3+4��f`X(9>7�U\�O!x�a�g�8 ����if=F�X��?2}����p��p��q��8�AX�3}�8��Yke�����P2�/"���a���Ef�ɬ�2���w2�C�X8;�C���xSƛ2ޔY�e�)3B0��a��EdXb����0�fx��0��?������q���q�����B�xQ����Q�/��G���A�� F�?
�B��(��
}���}���A�~X�.�<1���Q⛷��A��(����5�?*sSe}X��*Wyn��k�
g�s�
�ʬi0,ԇ5$��{p�����¹x��=��[�nH���ݕ#4�Qy���+� �°P2��pT榊�B,G��ƣu��*�T��p�0K,����s8 ��a�\�N�^�i��s8�ƣ0��w��x��X�B>W�|�X�6�ӆ��K�t���/8���h����p@>�Gc���8`!ȇa���J舣����lx%ð�+f=���1��9'>x�PT�q�M'3��p�x����+ꃧ����:��SN���8Yg�9p�¹�� ����:��N<�d&:�g��7��B���8N<�′8Nf��:y�:Y���zPG�/:1���t�љ��%�%ޝ�J��q���Wg���E� ��_tVh�tİ�+�3���0,ԙwݰ�¹諝>��cp\�3p�� G�O.�U����d,-Zb����GK\�$���B9qO�����a����!A$��>@B Ag�cx�H��O�B���Ez�H	� �W���*�E�H� 	-�!������@�H� 	`X����@"�?,�\� 	����g���q>A��+!�%^;�A�4H�$H�3�`�i����i�sAB� �W��
��ֈ먴�US�4�=��
	-���US��ܔ`�A�=H�i��U�=΅W���PBj��=�q	����4BB� �4B:�/���:AB� �=@�aH�	��� �*� ҁ���AB� �E� �	u����Pg|�`�B� A,$�����z	>!�'$4z	u�t������4B�FH��Z)��	���PH($����PH($(�3��H0)1ˠ3� �@Bg`X�+4�!��"H�U�	f %�<�@Bg %��e<��Pk����	 �!���'b�)�É�'� <���+�è��܄�@BC �$4\ABC`X8k-H�!� <@b_�H������	f �O��O��OD�Q�D�>�C?�O��1��Y۰�?�O��������!��س�
cxaED�?�?O!֟�����=�������}���"֟��'b��8~b?~"����׎_�<;�;�;�Q�������T��B&���5�������J�Hz"������T��h{"ڞ���J�'n>,���l���)��1�T���_yR &��k��w'�݉xw����^Y�TV�Ξ�Ğ�T�*k��}���)���]��BY�%OD�S�w*�C$=U�H�'��D�=[O($�%��DD>mΎO����D�|X�uf�!�3{�;�;�SÛ��XG5��w'�݉xw"ޝ�w'��'"��x"��w'�݉������}������8��(yB 7�$����'"鉸yB %OD���q�D�<�~E�'r=,�*�*��ľ�t�#����N|�x��p��N�$bىXv:��9���	}��>@"N�N�<� ��uB ��?��?���>��Lt;�NĲ��>@B ��X�e'bىXv�<_�N��ڇg��������ϝ��N'>,�Õ�牉'��'��(yb?~�������O��;���a�\q���3��Ll=[ϯbΨ�g������{f���X�WM��}&j�����LD>mϨ�gb������L�=[�5�����gv�gv�gv�gv�gb��}&F?,�+��2��3�aẢ�u�~�Q��D�3Q�L�>��?��)��Ld?����3q�LD>��xD�3��3��3����l�h{f?~&����g��yǛ�����3��3��L$=�󟉤g"陘xf�}&&��� ��1�L<�g?��Q�������g��3��~�Lt;��D�3����L�;����g��烙�(yfFW?�Eg�}f���p��đ��g��31�̞�L�<%�D�3Q�L�<%�D�3Q��.�L�<��Q������,�b��І�ygX8;����e42� �W�U�����pvf+����}FU ��d�D�3�U�L�>�*0,��E �A ��S|��2<@FU 'V��  �*�!��s1��� CdT2\A�+�(d��3�Q��&��&�(d��a��̰hdH��:AF� �N��24B�F���a� �AF� �!�� gV�0baXb}2�����lՐ�2��!gfs�Ða2��aX�!��ZB�a�0�aX�Ða2J�!�{��=�d4��dX���AF� �r�Q'Ȑ�!C>d2�7�W��+Ȱ�:"C>䂧�Bdȇ���=Ȱ�BɬrOv߁���݃��A�|�d+��&j��%��B�����a���
�J݃��A����"��`X��Lx���A�������^A���0�"CPdx�/�Q'��^"�Kd��Q�d+���l^"�*�!(��:�q�8΅Abd������"�!�<�Q�(���52�F��ȐcXhև�dT2DG��΅�Bkdh����52��"CYd����A���0�"��!CYd(���AF� ��!�i�a32$FF� ��!�W�Q'�hd�2d�	�����(d��ё!:�����(!g��2$C�dȐ���>2�GF� ��!Ádr@dȐLV�+�aE2Y!2�Hn�;�G��������#��aXbk����O�p $��!C�K�v42�
z$����F�h#d�a��I2<I���#z$��0,\�O�QT�d��d���J.eX8;���QT�(*d�/C�d2�,2�
R%C�d2YK�!y+24KF�!�Ր�j�/�%�Ր�[24K&�E�o���/��fX� �E���00�%C�d2Y��p�8�Vd2Pd���
D�o�(<d�K�b��f��,�ߒ�[24K�f��Bdt!24K�])d�(�,�R�4,'�W�*��]�@����R�Y
4KAq��8Q�[
|˰P�83���E�x)�K-��3,\i�+˫8W�+
�LA���\Q�k
���@�����E��)�T�G��NE��)P1�b9�O��N��wQ�d
�L��)p2��r�@��,
ZN���)�K!oE��);^	S�b�%�}�'SЗ(�(p2��*�@�2Y8�Bn�Bn���İPg|����8�Bފa�����Q�8��$
tM!#FAq�@���3,�>��*Ű�{�S�vQ`i
�̰�+��)��o:��Р(d�(09�����S`r
LNAˢ��x�oS�m
y4��L'SP�(hGș��D��)00�����a��x
|KA��@����RP�(00�\����SP��x�P1*�@�2k2kșa��x.�L��)00��S``��k��Y��k����(�+v��5�@�ؕ�RP�(�+����葂�E�')d�((`x��&F�0)oB7�@�(��R�P
�I!�F�9)0'����5�����P�(p)
���Q�P
J!GA[������R��(p).������R�R
\ʰpv<.����G�])�+R���Q`N
�I�����)&��a�5D��@�(��R`N
�IA�������@�����%�>�K)�$z�@�2b���*�A�I
J���8�BF���F!GF!GF!GF�0)d�(0'�<��P(��.���2b����G�')�$�l�l���L�����TK�v�7
<I�')�#z�@��=RP�(�9�Ʒ�V�@}���FG��(0E��Q�>
9)��r�����F��(��,݌�&F��(�]2Px�1 Qc/��%^tD!�CAˢ�K���s�3a*
�DA���1,��\ AQ (
E��(�:��BT2
*^bX�
����D��(�^��Kx��nFA7���Q��(�fT2

���\�����QP�Jf.�j(�(�(d�(���U0���,
\A�+(�e(�e('��3P��P�
AAݢ@�-
�
z�¹x�>y�FK$�C�F(��K�F(�Ҡ@�4
�A�=(�m�{P�Q�
�#��s���O(���qhtrRrR�K���0,\;��(r���"ǰ�bx.C!oEA����bX(����pՎ�P�
|BAmcX���Ρ�0K�R�XΉ�GK��a����*:�
�0�(9�+����0T�
�P!*�b��5���k�
�P�*|B�O��e�
�P�*|BE룒G���Q�*4BEmcX�W�~��
30,�*�h�B����T���F���f%�_俨P�l��a�>q�����B5�wȈQ�*4B�=�p����݉�WE����Q�*�-*\AEI��]��K��T����%�_��W"��\��~%�_��W������J�����=�<�<�B�1�W��Wb���J��%�G|+[ѩ�D�+:��J���JQ��W�9��h��EEˢ�e1,�=>�Tb��}%F_�Q��W"�|%�>,�^m�D�+�a�וb�����+1�DE_�%�䛨��+�%���Y�&Q��W�$*j�h{EM��&Q��W�$*��J�J��[�(ETb��z%�^�|�h>T2PT4*�����zC%�>,�P�aED�}Xb�"�^�[Q��W4*���Y5ef"�_T����}%�^��W��]�J�}X�R��l�B�x%1��Rİ�� q�a������Wb��zE�aXhU|��{%�^��Wt!*Y3*���
İ�b<��1,��%�ư����D�+�JD���D�+��B�x
�͇Jl���P��5d�B��QQ��D�+*�B9<w����d��h>T4*q��
DE�aX8^@d��5�ٯ��+��.D%"_Qo�D�+��zC%n^��W�*Z�ҟQ]�䭨�0�E�E��I�d����UeT'�^��W�]T�]W�:
ՅZ�Ϩ%T��(y%J>,ԇuJ�Hz%�^���?W�3�	��|%"_��W*1�J��JԾ��D�+�
m���*q�����Pg�y"���~%�_��g��݃J��{P��W"���Ps�-*1���A%�>,�!ބ�A%F_��Wb��h{%�^Q'�o"�^��W�	*���^A%�^�IQ�4�xD�+Q���AE����$�?,\�1b��X��PC|��%�_Q9��TT���`=E0,��+�����G�B#Th���A%�F�X�����
�P�*C%GEӠBT��
EP�*AEӠ����T(���A%gG%CG�+�p���`P�*��a��ޙ��������%�_��5�=@g��x�@%gG��� ��J�����pv�	���飒ţ�T��a��	���BE	���BTH�
WP�F�h#42}4H��ZB�=���FK��W���� J%�F��3�^���WЈ�7���,�U����A�h�4t\A�+hp���4��W��
\ACӠA4r4(�F����AC���`��
�>�A#�GC���W�`�>4B�=h�u�F�a�W�� Y<�A�4h�Ҡ��2�@���Pr�+��r�ە���=ʉ3c#?Ȱp�q�l�	>�����4BC�����=�W�݃�0,�9Ε�¹���F�a�<������Pw0A>4�
����`!�@
��NР#tD��h(4��4
�F��wѠ,ځ��`0,�OA堡r��7�F#�H��h�6�Ab4�J�B��،���Oh�%4�4(��6B��hp��F^�w1,�d��s��$ʢAY4�F��F����@��h����@>4tTC#GF#GF�shh�ħ���@�jʡ��ɢ�948��A#�Űp��ֱ�E��"hd�h(4X���@CC��04��� �BCC���L�%�D�+hP�B����?,��8���������ƾ�{�سߠA�h��oP�B���5R���]�����4��Kl��3��{�����a�\��W#�C#�?,����/�g����
��³9���P}�� E�P���M�/Php�`X(��"hh44����4���rx�f#�İ�r`�%^�$�%��N���س�س�س�س�س��
{���A�h�nh��op����l�B��^��7��7v�7�)4��!����:�ހh��W��%����Sh�JhD���yy<����a#�߈�7�4x�F��5�$��o��o�AhD�;�;������F��o�o�oD���Fd��od+hD�;���FԾ�S�����o�oD���F��o��%��l��}#j��V�ء��_�ء߈���U�Q���Fn�FԾ�g�����oD��1�F���o��o��Q�Fv�Fܼo��oDɇ�;�Iodh��o��odh��o��o��o����%���y#;@c�~cg}cg}c�|#J�P��x��o��������a�m��C��o������1�Ʈ���Ft��Z�9�]�]��vc�|#�݈w7�4�4"�����}�xwc}#~�>�w��8�n�D�O�ڟ�?�w��?�5��d�����x�Ɏ���'1��IL�$~?�e犾s�>���}�$=,�=�Ή��I�DW�$*}���$*}�������$�|��q>�8�D��%��n����I��$R|�ت�|Ob�';�Ob���3��DoO��'��O�'��O��O"�'��a�J#�t�=���{�Nb�'Z��B�~�l�=ٷ~�=٥~�6�ˉ�!z{�=��%�����>0��)�D�D��d����I4�D�~X�R|�h�I4�$R<,�#b'����ɞ����ɞ����I��$R|���<������PC|���I��d_�I4�d�I��$R|���$R<,���h�p��;;���+���N��'��'��'瓈���"}��&���'{�Ov�hݟĠO����?�J�D�O��'��Ov���΅��g�d���P�`��\尊c��p.Vz��?���D�O���ĻO��'��'����It{X8;>�b��b��>�������I�$�}��ت��D���''{�O����K�v��'��O��'q���Pg���';�O��'{�O��'*�'��O��g���ɾ��}�'��Ob�'��'������PC��h�ɾ�����.�������I��d_��Ē�D��$j��?,���ľ�����]��,x�����'���������N����Y�8"�'q�����5����I��$F�p�0,���|���I��d��I��D��$F����T���O"�'{�O��g�����0,�ÜB��D�D�$"��X(�^�SP�?�8���u������V��8+}5�a�}x�Bg�Dg�Dg�Dg�d���p.�3Q����'q���'q��8�I�$�?,��D�O��O"�'{�Ov��D�Ov��ag��I�Xhz8����""��?ٳ��?,�����ύ���f�D��D�D3�d��Id�d��I��$��?��?,�̊��M��?��D�O��'Q������a��<��� ��?���D�Ov֟D�O"�'��Ob�'1�����Ov͟D�Ov����X�x��O���D�O"�'����'�������
���џ��Ob�'��Ob�'1����'��O��'{�O��ǅRf��'1�a�W���~��}Xb�w�<{ۇŒi1z8{�O��'��Ob�';Ї��0��j�چ��I�~tL��?�ڟ�d?���d?����O����|'�މ�w"�HzG����������������;:���|'�މ�w��w��w��wv�wv�wv�wv�wv�w���8~'j߉�wb�����|gWx'�މ�wv|w�ww2�w"�Hzg�v'��э�h�w�nwvjw�e%���P�٩�٩��Y߉�w����۝8��P��41,�'��:<@G~X8{�S:��;��;:��}��`X�O�w:�����N�w:�@���
�0���sS�"�(���D3X(9�M���}��L�4�(�w(���W0,������h�w���X'�}'���9މ�w"��]ᝈ|'"߉�w��h{G!X�}���[���;
��}ٝ}ٝ=���Nl�I���;Q�N��%�����w��=�Nܼ%�(�w��w��(y'�|Gi��㻓k��㻳�m����߇��)D�;q�������P���N$��k�I��w��wb�Hzg�x'Jމ�w��;1�NL��d����;1�NL����w��(yGW�%�D�;�;*���f~gwyG�mJ���w��w��wb��Hz'Jމ�wt�;��;��N$�I���;q�Ξ�N$�I�D�;��;����~'��������٥>,��#&�Q���w����N$�7�Ǳ����߉�w��w"�����zGW�����A��]����N��ND�m���{�I�=��z'�މ�wb���Ύ�Ύ�N$���߉�wb�]�N$������މ�wt�;����y'J��k߉�w��w"靼���zg���ĳm������v��v��w������zGW��۽m�D�;J��h{'n��#��#��P?,ԙY�Hzg�|G��Wfb띝��h{g���+�"��B���C������׾���h�wt�;���{&q����a���xn"�߉�K�
�;<@��� ����{�������������;��;��a��Yױ�X80,���f��t������������������B�J��}���&b��}��8~g_g_'��Q�����D�;��N����D�;;�;��Nd��J���;<@gg�~��B`Xhy��]���wP���Xg_g_���X������������0�B���`:�@G3X�_�D�����댲}'������zg.�y�������wx���}g�~G���t��w(�EС:A�"��%3�����
:j ���~�F����!�a:�AGC�Ct��3�a:�@G���t�����'ز�z#�����ɲ��v��~��ޘ�0�,&���|��NL�J���^,������g�^P���ט�W���zU�U�D��3V[�z�f��e��봽N�zڙN�봪���w[�{��5���E��D�o���D{�������"XL4ή��!��� ���F�`1Y��}�u�]O���7<�b�(���*���Q9xc�����F������v�-�K��u�7��ɻ��a��ü��_LV©�Їވ#,&j85NM�s�0��excr;t�7��b�Ns��x8�z��v�C�Sӡ�С��(XL�����p�:t�C�y�N,&/�	�=���}�͆�Eg�7�ɖp�;�����1鏇�x菇��F�~1Q��̗t������xc�����&���@�b��&]4�����cr2L�hr~Lzmr2L:rґ��Τo'};��|�t,&;@�xg��#��-�M��&]4�V�5fҭ���/&�r�K�B�Gg�wo4��F#`1�C;yv����7��b����b+�s�='�s�+��D�4xcr��v�l���
��=�������*; g�(�rv�͎���˹f*��ѷ�1�]�8 G��ZD��8���b_->�����C���� �b��o����z��)��EM�GG�b�..W�˕���`P����W�o��ca�Q��1�cauM^�rձ���3rux���j/������P[�ʫ�ou*��.�.ӫݷ�}�r�GW�~�ct��W{t�GW� �5@��W��eAu$�.����S])T_=U���5yuV��U��9�7�������5���؜(�+��2����餹Lo�0Mwo�gj:r�k�^��ڦ�6W�MmN:M�m>I7���M�k��m>I7HMl�c��k��n����\�7]���٪9[5]��͵\s-����Z��p;���'�SG>u�SO;���)���N���U�����\{:מ.�N]�t�=��S<���Y��EO����t]x��;����S=u��uᩋ�N��o�O��S�=��S<�O����󩋞΢�.zꏧ��?��c�����%l���؝X�kwb�>nu}����W]��N�]G�΢]��cw��c����i݇��?v��;�vW��%l�k�^����ڷ��]G�>�u��o1�#@�ݻ�ޝ���ow� ]G�ε]G�:r�pd&��h����FM�������u�?������]�a]��a5YU��]ta7�_񰸿��vq�]�`>yj��.��K �����dY����~�@�_��w��9gj�Dw9���0�Je	%�B	��i�vV����.�0��x=MNa�SEY<���d������.������4��)컞��8�E��'�a�D����}�kv�}�Eо3?�2���3?����;O��dľ;������LM�d�.�KF��dU�����ud1��p;��C�=�Za��`���|���.�K3�3���0yA����<��(���d�~赇^+1L���:���0Y�ӯ��.��A��e��������C�9t���]�a]�E�C�J����.��'}(�0I�H��v��=9�%Fa7��vq�=�V��dYNM�e�inOz�l�����>�x�ۓ>���D��&��''0i��v��y(�E���%'���t>i�=�|�e��Þ]cf���K�=�T�y�3q�]�a��F��]�a�h��Z.;�HF�{v��؅%va�=�CY��z���.e��O�w{��3���0yAN:�I'�c�سxY��سXv�zZv]�]
��Y��:���.ױg+����iŇ2Q�������V�ӊs�@�0yFʊ�\ѷ�F��K�a����3_ѷ%I��"���EG.�|�&���^���M���8}[*e/:���^tѢ�]��Fe/�Pq]X\V��	L*e���T�.��W;y�y���eW�J�l�]�Uv�]e��{��:�U]Ae�.�� ����*�����9����T�.��K�앗��T�.�����UW�N:��D�d�z�$��`�vI�]�d�$�%IvI�]�c���˻f���E=vQ�]�co�����\�	q�g��b��,����^�\Y5�N�8v��]bcov_�����j��/v)�]�b?]F�.�Nߥ���d1vY���N]������.�1L�йC�b��O��e�,�~�C�>t:�Hl���t"�1L���te%ı����s�NA�c���E=�ӧ&��]<c��O�Y�]c���e1vY��$�;L6�K2Y��돲�,��}Uם���C��,�.���b���C�w|��!�;�uׅ]��c����]�Il�g��G�c���%6v��]<c�.�$6v�]<c���3v�]<c��/��,*e��T�EYVU�`?T��X�C~b��5�p����f�!�q^���š��!xq�,1L�����8d1Y�C5�C5�C<�x�����a���bj:T�8$6��+�a����+V��xơ@ġ��!xqHYJ?J?�<����!,qK�ޱ�z<�~8�y8v�C~�����Wu��ġ�ñ3�������!,qKb�
��á\�!�p(�p(�p�.;��!�p��p��p�%;Tp8�i�CNa��*˻Ct�P�a��۬��cׇ�C��p8"�C��8���2�2�d��4a�CX�P�8x�&�?�O������!�0jj%��d��C͈a��u8�.*�p�����w���!,q�V*8b�ġ��!qHF������!,q��0LTU~b����@����Cb���ޡ�¡�¡��!q��p$}HX��8$#ɈC2b��F'ä[��p$����u����\JF�U�oD��),qK��dUu>Ɉ#�CjFjFjFjF٥���!eqHY����ԟ8�sZ�	,&+���C������Gv29B�� #rȈ�AA �&����#;(��qBF��N�YG��8$6��a�u��
q���*�qq���ő/|ۉU��Cq��8q�)S��(
�A�8(�z����dUuQ�����g�zJx��8׊gj��ơ�!�q�r�b����!eqЇ�š�ǡ��!�1L��g*�ʁ�YTb�(�}�s��"��!�1L�j��PM��:��IrH����V��PF�9T.9B���	�����j#�d�\z�Gխ�n%r�j�!�2%�d����:��J�0B������"�\ǡh�!�q�#r�#r4���Ԥ��!r�*��5�
!GӭT9T9$II���C�	L��$9��Uӭ$I�?��z�ʁ�%Gs�Q!�Pd��F�DPI��9)r�j�%�p�!\r�rțʁ"(G�p+�"(������0qF�C�8�ӤR��kT9T9dWuD���v�g9�9dWBA�C9�a����My�a��ud�Cl�P��9Ng��E�r �r ǩ�	�j�%ǩ�.%II�C��C�d�(^��C��.9�K�?y�C9�C9�C�A9�S�T�!�r��ʁR)G�EU9�ΧhȡBȡB�!�rH���*���!�rH�����uQ�C���N��%GwU�c�,�YTU�CU�C�A9DP���w�]�a�t��ĚT�H�(�X�a��'�>��IR�#	�Sl�$I��Hb#Il$�jd��l&�a�L`I��$\��K��V�	,)��M��!�T#I�$I�$�?�BɄ$I폤��0����eR�#��$�?�TJ�JI
}$��$A�$���R�TJR�#����R�JR�#I�$U=��ɴ%I�%��$q�dڒ�BHR$)���Q�dW�zIq�$Β�Y�8K2�HR�c�� ֘Iq�$��^��K��G��$��$\��K�pI�+I���8G�JIR)I*%��$e7��0�'�Hf2I�u$3�$A�d&�$����&����M�ɲX&%<��IP%��$)Α�R�JI*%�}$�}$I�$��$y�dƐ$\�T�H&&{�>�^G�JI�&IF$	�$��$��ӉC�@H2�GRc#��#��#)���K���;��H�$Iٍ$\�L�L��M��Il$��$56��ȸDz�I�����0���C�I�n$�$\�$I�Jɼ"ɼ"I%�����eJ�$IR)I*e�,�գ��0Q{ٕ$���R�T�0qA٩Il$���*I�$I��!I�$	�$�$#2<��ȢI�#�z$Q�$ꑔIfXI!�d{���$EC�pI.IfkI���rPTIf~&+�JT�$���M��xk�\�B�0Y{G q�$ΒdW��f��J2�L�]&�(�2LTBv%)f�3Ij�$5I�$�$5I�e�,ޡCM�d*�$��$IB/I�%)-�dW��!���pPgI��}Bw/��8�0ل��
!�d%�~�I�+Iv%ɮ$A�a�:��$I�%��$��$	�a��
�$�L���0Y���&�Ir0I�%��2L��\kn�d"���IzIB/I1�$ᒤR�TJR�$�O'I�$�K��t��%�d%�Eͺ�* g2��0Y��f�L��s�L2yN2y�0Y�Χ��0QU9��
Jg&��8�0Y	�X%\���u+	�a����s�"+I&)��$\�9p�9p�ɲ��Dc�"+I&�)'����;�5=�����I25I�&I�$ј��J�I�1I&�)'��$јd�$�Dcҩ�ΒTgI�2IZ&)ؒh�>�V�%��$ٕ$���]I�*I���VJR+%��$q�$Β�<&�"PPe����p�
J�$q�a�}sj��$��dW��JR%���dW�Ij��J�]I"(Il$I$Q�d2�$�D=�������0IM�$���:�\GRZd�.ʲ%�;��RL,� IJ�$��$�E��G�HIb#Il$�$��I�Iѐ$���֒�Ò%6�xF�ȯXYeB��FV!$��_��&+��)�bp�fk&/��UV�#q�׈+�W��h�0Y<#�0Y�>qds�d�d��,ב&�Ǉ�:"Y�#��%�ud��lN���H��Ȣ�d%�!��d��a��&]��duD�xF���Y#^�]���"Yѐ��?L���&�1Lx�$�<,YM��3�dQ�l�,�3��a��a�!Y $�o��?��'Y�#�zdQ�l��,�1L�4�V $����?��GV�$��Y�#�zdQ�,�E=�:"Y�#�zd!�a�	�Ò%6��!Y#�a%�gd3�d3�d!�� I��&Z��ȇ� ���&J&��~/ב�:��"Yi�,���?�j#Y�#�ud�F�j#���#��Ɋ�d��a��ʁd�lҕ,���?�IW�@�0yF��ɥ��H��j�d���LIV�$�d��,6�U.ɒ$��/Y��,\�%I��$Y�$�d5I��HV�$���e��r��,Y�a���d���BH��ȂY포�G���
}d�,��M��%6��F���Yb#Kl��ҭT�Ȫzd!���GV�#�zdQ�,��:�9]�\G���rY�#^d��,e��֒�,��Y�"^d�@���l-�l-Y#�bd��,?��'�r ٜ.YX"Kda�,1LTB	�lj���G�y�Jx��ׇ��IW�IW���0Y�>d���^G�Ȋsd�l��,����R�z�d��
bYb�.��ui�,�����S��Y!K ��@�Y!��1LVB��i�Y��,�����Y��,�0L�Q��f�Jxd�:�zY���^G�yȊsdх�G�S�*qdхa�>��.dS�dU=��CV�#�<d����G6�KV$+����4CV�c��jӷM�%#�i^�dD�����\�I3di�,͐����YU�a�*��� ��C�f�
}d�a�x���|Y�!8d�,͐MR3L�4'�U�f��M�U4$KFdB�dD��bٌ4Y�!�<di�,͐��4CV�#������bY9�a��ε��d�2�[3L�Q��Ȓ��2�d�\c*��U��"Y�"�E&+�1L6�nu:
Kd�>��e��Y~"�X&Kd�>��e�HE������2Y��a�x)���GV�#^de7��EVv#��%��%��%^d�2�������<,Y]�a�@P#�Oda��zF��&/ȥ��Y��3�
�g+u1��E�Ȃ��
��l-Y#�b��pj��(&�)B�d0E�����u!�"�QL�R��(BE�c�,O+r�d0E	�b��"�QT�(��a��E����QD=�JE��H鏢^G1eL1eL)!��2EFd���^T)�$�\3E9�b��"RB�@H1#�0�^�)
}U=�@HQ����Q�F��H)�)�$�d%xS�K����5��;����GQ裘ʦH���"�R�R���0٪"(Eޤ�ᒢHQ�c�l/�j׭D=�����m�l/݊��0Y	��@H1�M1�M�)*���b"6R�[SLRS$I�$I�$)�$E��(R)*�B��l�Ij��IQ�H���"#RdD�i��El���Q�L�a�Y��a�,�O�țy�"oR�M��J�|J��"�2L���oQm�țy�a���&Eޤ�IR���LI1��0Y	F�����ҭ�K�pI)
���"6RdD��H1�M)f�)�$E��a�}%I�2%E��b�r�0��}�R��&��9��9Ev��)�(fRdW��$EM�b�"�R�))r0�DYr0E��a�q̧3L\��L��)�2�dY��TJA)f�)"(E�bb�a�u>�@�$I�$)�9M����GQ�(�Q�K��E	�b��a����$EF�(�Q��(�nS���"6RB�i^���0qFu1���D�T�(�<,E��bҕ"�Q̰2L���ư\�� ��b�t*Ebc�<�]���Rˢ�u!���E��(rEŋ��E�(
WT�ղ(jY�+�yX��H�&j/6R�F��H�)2"EF�Ȉ�-��H1�K)b#EF���ר#�楈���#6R��(Je��"#2L���;��.6R�F�"E����!���EQ���RQ��&�Q�:��FQ�b����F��(�T��'�\�i�F���E��(R�d%|Ql��a��,QT�(R���`�D1��0Y��!�)�",QԌ&��YA~�K�g�T�(*Kө5#��E��(�S)�E~��Oa�b:�b�"R1LV�IG�^U*��:QHY)���D�("EX�K�'�ɖ�QD����D��&[BO;��'��D9�Ѣ�DY��DCw���C1�Hp(�He$�4�0Y���$"Ee���D1��X�Z�=Z����D1�HQ��(#QD*����9�HYa�"Q$#J���}d�� ��,��E�b�l�N� �Dp(&)2U���.TU*�)?LO�f�bKT�-�)^c5mI5GI5GI5GI����UX�
KTa��F������q�a�h�����L&�L&U~�JFTu1�Dp��U���.T/��N��Uy�*�PM[Rղ�jYT3�T�-��Cp��`T��TӖT��a�^�UN�
%T��j����EJ�B	U(�
%T�3��[+�Pw}H]�*�P%��0Y<1�*�PU���;��`��ȔY�&��*�Q���@��UX�*�Q�'��D���@&�%�0L��p���RUj��RQU��R�D{�}��eQ�>R%��^(�0LVBO]�B	Մ$�Ї'09�*�P���B�S�r
����3��N��BJ�B	U(��Tq�a�^z����*�P�Ũ�bT�-��0Q/q��\=J Tu1��U]�j���.F�S�JeTх*�P���|'U��
Ԥ�Tق*[Pe�lA��F��bհ~5�_M[R�פØ��ï�坩F��j���&.ȼ"�P|5�H5:_���F�a�%T���HTc���0�ɳ�\e�j���*K�M�+(#Q���re�f�0Y�s���jX���s�bUe���D5�_M�Q��QU��RU�jJ�*HP	��U��*6Q����&Z�,U(�*IQ��Q��1L\c�8�I3Ԣo�xQU�������bTӃTT�2�HEU�JYT)�a�x�ӊ��U]�jƐ*x1L�堠TF5=H�UA�*�Q�8���0�8N�BUٍ*�QM"R/��E�&k�Px�Y��-�QU���U��*�Q��BU���jd��FY�*�Qe1��rq*�1L���G%<�xF����U~�*�QE*��D5c�0Y{]T���TT�8�H�0�8��U���zFU=�*�Q�,��A��,�*x1L����dYN��U�
^TӃר�F�Ũ�Uٍa�z�GUv���Q�ب�ռ"U�ctBk�̧zF���BU��
qT���.FU�
qT!��TF5=HU��zT��*�Q�ŨrU��*�Q�ʨJeT���TF��rU��
qTE0��A��0yFO�8���|��JeT���zF����dUu>S�TQ�a�Ns�.z����#U �JTQ���FU*��uT��g�;N�&�-�@H&:@��KT�a�,Wi2"Uŋ*6R�F��3:[	����<$\R�Q2L���T��*6R�F�9J�9J�pI.��uT�*\R��&7�*qT�*\R%I��ڻ.�*qT�8�J�d��7��&Uٍ��F�J�R)MޤI�4���z�0�365��HSc�)�ф8��J��kBMb�����)��L�Ҥ?��GS*c�<#>Ԕ�h!M �)�є���oY/^m6Q�fr�&��Բh�M�c�,��\�hB�D%�:�\GSˢ�u�-�ф8��M���b4Y��@D��h�M��&��L5�/��E�h"M���j�IY4)�a��;��E��hJR4�4�'�H�0yF桦$ES��?��3���d{153�4����D�&�7�IS���R�T�h�T4�&I��F��Ml���4��a�,�9�fV�f
�f��a����o�M���z4Q�&��D=��kd��D=��G3wJ��h
W�7M�3Ji��dU�G%)��H�i2"M�a�U�&ΨpES��I���[�a�q��&#�D=�*�(�(M�a�(�r5�ISˢ�e��h�%M��I�4I�&I�$I��M�d����&o��M��ISF�����4���DSl�I�4���D�J&����|gi�,M�&�Ҳs�2Mve�����0Y�3��T��KS��I�4	�f�&�2L^��,�Dc�IW�hLS�I�4u1�IW�Ɇ��U�h�g4�4����FSc���4��f���FSc��ӥ	�4a�a���7�.M̦�����4�:� MSv�I�4i�a��fki�1M�	�4%<�L3�K�iũ\Z�I�4јa�^N��4��&���Y��!�4/M��&��U�9]��JTiJ�4�4U=��HS����4��a�,�GI�&I�$I�$IS��)�фK�pI.i�%M���X�	�4�@�B��0M����43�4�>��Hi�tiJx4%<ZuU[���h�&��/M�����U��$�d{53��gtjAi"(�d�\ժ��DP�JS�c����h�&o�L����2L���G.ij4��ݜ��R�TJ�J���l	���t&��ɛ�Uu]h��fj�&6�i��4EC��I35K35K�JiR)Mޤɛ4�f��%�˙O�ɛ4EC�pIS4�I����pIS!��t�	�4�f�&\҄K�pI.i�%M��a�	O����e;�I�4�a�x)�R�T��%6��GA��&IS����	�4��&����2L^���b&M�e�<����K�pi��4S�4�M��&t�0�L���Z{W�&�i&�i&�&[���\3��V�I�4�X��fZw�P����4��&���s��&4oM��iR<M��)�2L��@��45\��M�i25M������]i�2��6M�f�p5\�R,�T6M���ݦ�Դ����4i�fޚ&ӄ^����i����3�/�4�̩:˩��0]|�z��Oi�a�̢�"+�"+�"+��*�0�0Y/Vȧ��0śv*�rJ�J����9e}N��S�g�l/&�S���9e}N�_N��&�9�[s*�r�~��9{N)�S���9M,s��
��
���=�IjN5\N5\N�Ӽ5��Ϲ3?��?�ykN�S�g��_��9����3�ۊ��rC���)$t
	�&�&륧		�J��BB��й�y��rJ�R<�Z)�Z)�Z)�Z)���)�3L�Q��Y���7�)cN�Ü�8�D%�qNa�Sg���0�)�s
���rU��9ՃO�V�5�D�i��S�g���.�j�)�s*�r*�r*�r:�ykN�ԜA�1�d���J���;���rC��Щj�iS��4�)7t��rC��e;N�@s�@s�@s�%�bI��rNujNI�S,�K:e�N�S��4yΩ(ͩ�iӄ7��ѩNͩNͩN�)�t�%��r�^:թ9��N��|:�7�<�)�t�3���9��9%�N�a��ĒN��S,i�<��nZ�S��Sx�T�A&[BM�hr�-�tJ*���9́s�3��L���)�tJ*��J��rN3�j��L�Z<�Z<���0q�&�&Ϩ#g'|y�SŞa���J���)�tJ*�����K���0���Ny�S��T��^:U�9U�9%�N�N�NI�SR�8::�N����r8&�r�U��T��.:��N�wN�S�a�(�;$Jt���D�b9�28���Y�G�qN��gtb-.��N��S��TR�A:��9ŒN����F�*;���)�t*�3L^��X����yA�S�T��T��4U�)5L^�3��NUv�ɖp��:ťNq�S�TR�z:��N�S�i�pd��S��S�Te甍:�9�9%�N	���I��<��;��;�թ��)Tu�K�f<:%�N	�ӼH�d%��9�N�~N�~��z�LW���:�NA�ӌGgu��:�NA�a���E��9e�N�wN� ��P�Z<� �)uJ=���M��:͞t�=�T��z&���(u�F�j��&T:U�9U�9ťNq�S\j�,�	L\��&+�[5g>�.���T���|�$Tu
U�T�d�j��N��a�	udѫS��4_�)Tu
U��]:��N�.��]:%�N�yN��S�j����aq�S\��:��9%���p��rV���)gu�Y�
�
��r��:�:��NѫӤQ��]!�^��W���).u�K����%���z�h>���N��S�ꔠ:ťNq�a��ʅ�N��N��S��q:E�N�S��g&n�BE��D�)�N��F�Z	�]6�T���:ťNq�S��a�:rw��m9�a�:��E��E���)�uJc��X��e�RP�4�֩�)�u*�tJv���:%�NɮSi�a��
�^�ٹN��S�S$��bYЅ��ٹ��W���&��j*u��n����R#����EºHX7�V���]]��Kvu���W�&o�tWy��^ue��4V���j*u����0yF����\]}�n®.����Օl&�gv�"a��52�w)���S7�WW���u��.8�Ǻ"Q}�-YW���u埆����dW���&��&�&kϲ�K�uե�2Ǫ:(Ȓu��u�a��'�����T]�l��l�	e��xYWp�+8ՅкRR]�����˺xY/�JIu���ZWJ���k�<#oܺ�Q��_]z��u!�a��!�%�օк�Y�8�g]����uY�.K�eɺ�X��JIw[���[�+%Օ�&/H5�X�%�0�?ʒu5���>�T�RU�8�Wu!�.q�%κ�T]Y�.q6L��qB������@�o+^�Eº�U]$��T�EºH�0yF'ie���T]Y�.^�U��&8�g]p��g�eɺ�X�c�4h�4h�dK8�H�u��a��N�Bh]�K�u����VWA����+�Փ�
Z]�.��EՆ�r�H
ri].��u��rY�tQ��Ń
Z]m�,�	?9��u��a�Y�Vk��F)�.%�EºHX7�[��
au�����u+���VW���u��.�Eº�W7�[W��+^Յ��JU]ث{�gt�V��Kvu��n�nz�.����֕��fl�Ku��.��U���_��l]$���u���YֺYֆɲ\Z�A�Ǻ�XW7���M�֕��c]��Kvu�ua�n�.��e���kt���b\]f��lu�.�ե���T�d{���b\]��hu�.�����W]f��lu�u���xUW���lu����U��&�&�M]�ՠ�RO]�K=u�.�ԅ��XR7�XK�*Bu�u����N]���3uy�n��^]l���K=�g��+5L���P��$���̺�R]Ϊ�Yu9�.g��y֕��W]��nf��xU����X��h������4V����O�Wu��.��͌�Ÿ��V��Z]=�n��n��a��vɮ.�5L��գ�W]���qu����Uo0�b�b\]f�hui�a���q�,k]���x�+��e���V7[��*huɮa��ju3�us�ua��\V��Wu�nJ�.gՅ���S7�Y^�J���!�.��Œ�ɖ�;Nׅ�Du�.��噺<S^�Du��n��.]4Lԫ�}M��Œ�ZO]�����0q�z�"N]�i��l���>S�g�bI],����͟�%���N]R�K*���%���0yF�Q,��x�K*uI�.�4L�mg>�.�ԅ���R�T�J]R�K*uI�.��%���T]x�+K�噆ɪ:�J=uū�9��z�&7�[7�[�z�RO���WӴk:4ULqʜ&G�i*��jM�)k�^q9<Lq��&����4Y|�������1g��Ds��z�1g��W`�ɖ�c�4Y�8�S:����`��}��&���4YVt�a�˂i�����dKD����&ˊ�<Me�:2�W���z5Mt&��i�^PO�d�qY0L�Qw�hUx�i���,�&/[��c8e��0H�_cM���e�4yAz-��4yٺ(��4Y�8�O���ᙦ���=M�W����J�ȀP�d��<Lz-<�4y���;L:2��4y�q��&�J��i�	����C=M�gt���&j��X��uw�i�x�m@�i�H�7M�ީ�i���o#�5L�ȀP�d��u�09�"q5M^���4L:2�W�dY�#zV�d�N��YM����4M���%M�x�4Qդׂ%MM�4L���.���4Y�.
�4M�X�4Y{]�h�,^�E�j�,�E3�U�d��pC�dU�~Q��&+�#�z5L.�S|�&��ݓ�Mʾi����4yFG �a�ݡ����ѷQ�&�� Ri��i.����&~�4M\��4]��k$?�4�-�6�`Iä�M��,���4YU��`I�d%�k���&+_����4M��ji��&zmv�F�j�������4yF��d�&�m���ɛ�o�o�l��k��*��4Q<�U�D��YM�
�4M44��09?�G4�����|`I��{&���ɲ���}xi�l	}��i��|�DM�ר[!�4M^��P�ӊ�A�i���U�4Y/'Cx�aҭ�����a��������J %5M�RR�d���&�w	���4Y�3_u%���4Y��HN�i���AB�i��i�#�N�dK�8�&���ٛ&륧�YM����8M�ŷ�_���4y�>�5g�����A���3�o�,�<P�i�:�O�dYzG�;������A����$��&h�F�i����?�dU�р=�dY� %��4y;���l&�d�>���a���3�J��&��Ӡx��"�4Q<I���}��d�4q��>ä[��n�����d�4Y��BĘ��x�KG�.�&Ϩ�"�4M6���4M���&��&}M�i�x'0��M���
��I��%�K�t�C/H�Fyi�|o�4M��#�8M-A
�a�k�$7M��i�^.!���&K&�c�%M�e�0H�d�.a���3��F
�i�x���t�������5&��4y�z-��4Y/]�h����S��a�E����Iz7L����&[��<x�ϸ	�BB;�G�dYL��DЎ��4Y��	����&���Nһi������?���.س��R<�dY̵�`�.ų��n��=^���mϛ�]�gGi��l�vG�h�<#K�]Hh&����]HhڑF�&�����4LLһtю�4yFF�]�h�&�q��w�.ڥ�v���ar�@Si�<��	������T��g�&�1Gi8ڑF�&[���.���G��e;N��o�,�e�hz�b�&o3�.J���o�<#�ۻ��.p�#�4M��z��QK&y'J��D���.$��]4M��w g4Lz��0�8�=;BE�DC�]4M�,ųK��ƛ&��Э�3&gd��]�gG�h�,޹�<x�dUu>��]"h���p7LΏR<;D�d%�!R�M�g�a�J7MV�E�ѱ'׾HM�����9;JB�d%�t�&����sv���3�IEh��4�~���y��{���v-�'�V�gG�g�,���A�i�Uud��M�7�)��i�x�G��%�i�^N��=�`�.س��=��.ų��n�(�Du�DJ��";���N�i� �e'�B�d�|�Eoh�t�쌌*�4�����&��$-��6n���.*���4M���Sɛ]�f���7M��>$f�����M���i��S&�B���l���In��*�BäÈ��b6;�B�DK�$4M4N����&�茌��4Y	]��u�d%�G��]nh���v䌦�J8#��M���>zG�h�<�Ϣ�M��-��K�(M��;I#g4M��qB�h8&k�8���4�-���|s��		�BB���Nr�i�x}9�i�΢U%G�09e��rC���.7���rC;2Kä׊��,M�g�EQ^�&/HO�.�E���❤�v��a��(��ɩ��i��Z���I�E�i�<�>�N��]4W�ťv����J��F���%�v	�]\j��ɖ7L��l�&�w�G�i�h/Ę���i0�1�����0yFG$����v4��e���М���ɪ:o��o����bL��u����e�vi���z�dU�l�&+�-���fo����M��i�����c�&.H�k�8�d�.ٵ��o�twɮ]�k��&��8A~�i����"Q�d%\�H��Rb�H�.쵓So��� ���2[;RR�L1�ɞ� ��i�39(Hv�]�d��Ѫɪ:N���^+�����E�v2�M?��Q��&Zu�i��KM�]�#85M�G��]�k����v��M����v]�4{�d%tѮ�vgwY�]pl��cґ��&�7����4Y	}[fk���vT��ɲ�E�77M?���4��M��r�D�i��lK�2K��)�u�\n�.���8u]4�&<Tq:���&+��y�l
;b\��N��֡�ӡ��!�u�q�3b\s[�&��:�7wrV�P�!.u(�t�In����٨C6� ��4Y	<�g:�F:��M�gd2<���Cx�^:Ēu�I�CR�A:d����To�dYz�jI���i��e�fPG�-��CѣCR�A��I5Y�}�M�e��;d��C��P�� =�4Y<�2�M�g�EwV����!�t�pt��m�(�p�S��P�� c�4Q	y�CU��\l�B�*Tt�8"N��D��D�d%t>�Cx�^:��6M^��2�M�g��0yA<ROIܦ�z�dl�&��d(�tz-Y֦ɲ�Z���������C	�C	�C,�K:Ē�����m��lU���C��P��q:�y6M�RQ��g:䙆���G���e���G�Cq�C,�K:�S6����%�.&ט*	�����t�0٪N�2H�d�U6h�<#O���A�i�u��zUq�C�A��e9�� ���J�D�D�<�!�tH*�J���!�t�%��J���AJ�i�.t�.:*:��U�R�M�gtb%��4Y��aA�C	����n;��F�b&�Z%�٨��ksM�e��Q��D��D��D�D�T��!AuHP�BU�
G�P�!AuHPT�l�!uB�P�ئ���m2�M����[�Z�����Ci�C��^:���Cx�^:�T:TK:��Cxi�,�b��M����c:�Ř٨C6�P��P�� G�|�,'��8A���CYBU�P�0Q���!gu�Y�1d��&�wYP]Hc�X���!zu�^BU�D�Vfi�������!.u�K���$]Hg7L��l�A��i�x�rA�C}�C��:���C��P��g:����M�M��%�8���&�^:���C��C��CR�T:H7M4��N��A��i�x���tѡH�Aڸi�%t>E���J��K:Ē���u�uH*�J�d�d�&gdy�Cu�Cx�^:��2�M�e�@,]t�rC���0Q�(�A�����3:͑�m��CA�DС"ԡ��!t�n�l	�9Y�C��C��a���S��:ԍ:ԍ&��o��n���ӯ�S��S��S���!�t�E�tѡH�!]t(5L����冎ӇXQ�CɦC"h��l!�C"�&����!$t	��p�*t�u	�DrC�d�\�
	�KrC��С��!$t��n��m!�CHh�lU]T�� ��4�к(I��k�k�:��S��ҡ��A���xW�䛛&k���.u�8�K���!�tH*�JIE�$�����"QI�)�%%�dڸ$��d��+�6	S�9I�(I%Q�d&��nT8J�&����Ē�XR2m\Rpj����L�D��ɖ���TI�$�ԠJ�RI��U2+]��JrVI��$z��]�D��JUI+)K���J�R%��$��d��+��T����WR�*Iv%ɮ�xU2^R�*��%a�dһ$������S��xIu�$�5L��z"	{%a��,U�J��K��K�_I�+�%��d�$�D����d����U�%K�cIp,	����0�;��/)��LƗLƗDՒ�ZUK��KriI.-ɥ%��$���ҒZR+I����8�\V2�^UK�j$ЖL�7L���Z��]���%岒xYR.+I�%Y��6V/K�e�<xI�,����˒,Y�KRbI!�$%�����T~�V�dI��$K�L���˒x�0�u+u��:[I���VRA+	�%E��@[�KK��KriI�,I�%�d��$8�ǒrYI�,��.����˒rY�d%tQ!�$����J
a�e9?��.	�%!�$���Jg�d{9e����ҒWI-I�%��$��J�^I�+)K��7�D)���TI�a₲n%%��Ē�X�Ns�cIJ,I�%����X�KRbIJ,I�%)�$%�Lz��ĒI�I�,Y�K�e%��$8�ǒ�XK��K�dI�$^�Lz�$Β�Y�8KYw�8KgI�,�/�ٕ��J�jIT-��%5����0Y	�ʕ�J�x�-�`������Y2�^*>#��$q6L�K�TsT�J�jI�a�����JgI�,ɒ%Y��\�0Y��,8��ĒHX	K"aI�+�f/�q%��$��d��zV��xI�k�C<��Pt1�T��%��
Z��Ÿ�W�N�2[I��a򌺕dW��Jf�Kf�K�l%3�%ɮa�,�i$����VRk�,^�K�_�d|I$,��/)��ǒ�XK�cI5�$K�T�J�q%��V/K�eI��$q6L^��tu4�8&�w�PT+ɥ%E���XI!�$�6N�js}/���ВZBK�e%!�$��L8��.�DՒ�ZRT+��%岒ZR+��5L^�+w����Z2yaU&�ˡCz-I�%�a�̍�L���גY��ZBKBhI�,I�%U���YR+��0)���+d����Z2�a2�aR+	�%��$Ж�ג�WI=��xUUK�jI��$����J�R%�$�6L�Q�^K�jI.-	�%��$^�ǒ�XR�*ɒ%������r�V�*	�%U��\ZR�*I�%�&%��WIT-��p����-��T�d܆ɲ��OY.I�%I�$	���J�pI.)��$��z���K�qI�$/��咼\��K�e%I�dRŤ6VR+I��gtv�K*h%�*���y��IT-��%��$���Jf=L�8L�jI5�$��DՆ���8�@WhK�KL2nI���W��&+�С�W�K"t�<���3�b��xƬ�WV�++�E販��32tdA�l�Ƭ��0Y/VY����W6gc��&�g��&h�"t��Y�.��e��$X6Ac�˪�e����C���mY�-K�e鵬��0]�eU���0Y<+�,���Ҳ\Z�%�"aY���JX��3̂cYp,���g�U	˲dY�,8�˲dY�,˒�M�$�U�BhYű,q�eɲY�xY˂c�܈٬�YJ,�L�Y$,�eEȲ���b�|��d�|b\Y�+�qe��JX6ya��
�eɮ,�5L�^k�(^y�,�5L�Ţ9�leU��i&B�b\Y�+��U	˒]Y�+��0Kve��,����2[Yf+��p��_f=̒]Y�+�i�]Y�+�6LVB<XGg��,�E²dW���fP�fP�2[Yűl"Ĭ�X��
�Mh"Ĭ�WV�+�q��p���2[Y��,ƕŸ��aY�+he�,����f��,������`YI�,����&/�ZY��l��l��,ƕ�˒]��Y�+{e�Ų���bYy���X�%�ʋe�Ų�Y�8�gY�,+�ǲZbY-�,86LTU�,�e)�,%��ĲZbYp,�e��,8�ǲ�X�ٹV�++6L����܈Y�+{ea�,�ͳ������0yF�ɮl��,ƕe����0Y��I��V��Z�ԋYy�,��e���UVq,�8���
�e1�,ƕe��4V����XY�,��E��ZbY�*�%���fP�ʋe�*f�*fEȆ�z� 7�b6�bV�,�e�,f���.Y6�b�%�J�e�,^6L6����Y�8�ʋe�ŲZbY-�%���g����ͳ��g�DU%β�aY�,+��˲xY/��eY�,��1�e��a�
j�e�Ĳ,Y6gc˦^̦^��eY�,˒eǲ�cY�l����.q�%β�Y�8��eY�,��1K�e��,q�%β�Y/��qB�,+h�4�BhY-��1�e!�lfǬ�Y�8�*�e�8f�8fQ��^Z�^&n�jY�-���ڲ@[V/-��e�=�m��,���ײ�Z6��0Y{�Q���Z�K�riY.-˒eY�l��,K�Gˊ�e4f񲬄Z�8��l̲d�dU���˲,Y�%�
����eɲJhY�,�g1K�e��,q�%β�YV/-K��0Ac�K�QVBUh-�e�Ҳ\�0Y/�O-K�e%ԲxY/��eY�,+U�%βxY/��eY�,�T1K�e)�l��,%��Ć��2ǲ��0yAN��eY�,˒e�1f�1fU��Ӽ��݅в�kY-��1��1�e!�,��Uh�riY�,�e���Z6�b���*�e�вJhY$,Kve5βgY�+{e�˲Re��5��^Y�+{ea�,ƕM��%��W��Z�d%�!�,��E���dY�*U�ʆ)��(UVD���eE��^V���PU�*&U,BUE��HP���V�܈E��a�,��".U�� TQ^l�,�ɰ(/V�+ʋ�ĊZbE��(V+rVEΪU��`�,rVEΪ���aE���^�Æ�z��E��(	V��*�WEΪ�zq�8�PU�*
t	�"AU$��U��*TE�j�l	�Q��(�Uv�Y���PUQ����Uv�V��HP���:[Em�".U��*�e���\V��*rVEΪ�����:[E@�hi�bfǢ�V��G��"�Ud��
ZE��^�=�CG>���ѫb�Ǣ�V1��0yF�]fk����-�U��&륻{a�"�5LVBG6�c��*�q,�q&[U��*�^�tQ�wHw�*�]E���q����2[������*fv&�*zUD��
ZE���UL�X��Su���3�Xĸ�j\E��Hvɮ�@W�*�j�8�8��,jf�"�U��aa�"�U�Y$���[E�k���n��V��&륧Ic�7��P@�Hc��w24gc�*BUE�"g5L\��]�̎E@�h����V��*2[E@�(�U�.*AU$���z9�z�(�U�*rVEΪ�����Uĥ���v	�6V�*�R�d���R%���*�^٨��UQ�j����'�TD���T�ԋE��"�TL�X�� T�*�P����5�T�(�U���BXE!�"gU䬊zVE6�B��"�T䙊<SQ���3U��<S�g*�LEm�a�cJ*�e�-�cq�,.NE���S�g*�j3(�K��>,��U�J�k����R^*�KE��"�TL�X䙊<S1��ٞQ�S�� �����0Y��'�TT�*bIE,��%!I�"�T$��XRQ�� ū���0yA:�)�TE֧��Y�"�3L��h��"�S�*�?E�����"�SL�X���OQ�����a�^AE��"�S���O�&���(�S��������-�ST�*�=E)�"�S�*�=E>���S���PEdg���>$�S��|R<�d�Ns�=E��"�Sd}�RRE֧�����"�SDv��N��&+�f��a��{���PE��������$yS�XLX$o� M1�_��)�3���LM1�_�)b6E̦������󌺕 M��)�,��a�9������hL�)J6U�)r0E�(�T�T*
(���HEZ���T�e��L��)J#�3����Q������"SSL%X�8L�׊���ɛa���X�X�q�0N1I�0Y��SQf����e9?J�)���R�)�=EM�"�Sd}�`OU@�
�S�}U����T��*�SM8X�F�R<U��*�T�TX�F�J#U�V���:H��U֧��TM8XUK�AU���]���TY��ZR��
(U��*�Se}����JU�g�,w��?U����TY���R���?U���7��7���T�j���>S5�_5�_Uũ�U�������MU���UQ�*J4L���P�X�XŒ�XR8��EUɦ*pT���MU�
U�����bLU����TU^�&㫊1U�j��*74L��JU����Oݙ~�`O��R<U奪�R5�^U����T�U�U%����0Y/�V�*]4L���]��*pT���Q8��D�DH�
	U!��HT5�_%��DU���U3V����z�,P]�� Uե�XRK�bIUY�*�4LV���j��*]T����P��~�dU�X}�d|U�
��S�A�f�I�M���R�T���&�K���3Uy�a�^���RU��*�TŒ��SUu���T5o`^��JUR��%U5����0yAz��R5�`U��*^UE���UU꩚]�
BU����SUϪJ=U���JU59�+%U����LU��*�T%��	�	��⅗��R�T�bIU�� U�w[ݨa��.�噪<S�g�f��JUR���J*U3V�����"QU��*�T���S�T�&��&��j=U����RUũ�%U%���L5�ibIU,��%U����Z\�%U�Zt+��*�T���Q8�GUਚf���Tv�
;բ��4L6�ne2�*�T�T�bIU�
U5���JU,��4I�*�T�Y�2HU�� �g����RK��1UŘ�bLՌ�Ռ�Uɦa����z�ŉU�*�TM%Xe����lT����PU��J��FU٨ZMT��*BU�������OUa�j*�*zU嬪�UU�i�,�u��U��rVUΪ�YU9�*gU��rVUa���SUة*�T����M��])hU��U��*�Ue���V5I`�٪f�����WUΪ�YU9�*gU���U���&���쫊���x�Oѣ���0yA���T���Q�,~U�a�x_c5]��~U��
UUՒ�������JU@�Jc���Ӛpe�j���Y&�ީ\�k�<�S�����W�쪦���^U��*�TŸ��MUɦ�dS���]��Uث
{Ua�*�U�g�*/US	��Tnv�jv�*^V�˪�OU⬊��ӡC��a�,G���]��*�V�҆��}Ȑ^��k���T��d�:N�m�jv��nT5��0Y{�(�ު��0Y	gwu���[{�boU��*	W���pU�ʸU�VQ���S�^��jռ��$�U}�*�V�ЪZU���د��T��WEժ����Z�^��kU.�ʥU��j����.���DU�*�V�Ҫ\Z�K&��EMXڪ@[h��kU����T5I`�K�riU.�ʥU��*�V��W�jriM.�ɥ5ե�)�WSp�����A�L��L��$�$\{k2nMƭI�5Q��U3e_S��)K5LV��&���j�kMY�&���Қ\ZBkf�kriMu���T�KkriM�&�6L6���Қ\ZBkgM⬉��W�{S��	�5!�&�քКZ�8k�W5�6��&^�L�Գ&������Gū��UM��&K�dɚ,Yk�W���vS���믙�)K5L���&q��jfl�Y5����USϪ�g��ҚZSϪ�g5L6��,��Գ&k�#�z��TM��I�5Q��RUUk�jM�����2o`S��N��e�d�x	�T�j*U5���xY��j�l�_M���7�)8�$��d�0Y�.*�5L6��x8�
{55���S�$���Mث��L���Z��+%5L�K���q51�&�����䬚"QMΪ�Y5埚�U��j��k&�k�RM\j���
;5q�&.�d��l�0�ɓ�U��j�PMj�<�S��S�zjj=5A�&�L���j�D5��PU3��0Y�Os�i�&z�D���QM������k�j�XM��&��D���U��&���S�j��k��kZM@��.5L��AA��&��ĸ�W�jb\M�&�����T͔}M����T�j�^Mث	{5a��'L�ׄ���TM����gԷ忚�W��j��k�^MY��,U	k"a�D%D�W�jb\Mf�)%5L�m��5��dW��j&�k�R5e���������UMp�I�5)�&֔�j�_͜zMث�A�ԠjjP5a�V|�#��d���V+���V��jZ��]��l5��&���j2[M�&�դ��4V��jBUM��	U5e��PUS��IP5	�&A�ĥ��z���kTM��&�T�j�P�<xM6��F5٨�RU�j�QͤwM\�)^��]��]פ���S�z&��[Xū��UM\��g5LVU�f�&.��J�T�j�R5��a�f�k*U5���4VS���T�LT���4V��jBUͬtMΪ�Y59�&g��jrV��e���7�͇k��Zs�jZM@�	h����\��Y5��&T5L�K���j�RMꩩg�ԳjROM꩙���35�&��L�L7L��(�����Q3��0q;�7�d���0yF�Om�&�Ԕ�j����R�Tj2H��uM�f�&��Lg�Lg�T�j"NM���W�g��z�ε�q5���V3w]Kj&�k2H�Duͬt��-^ߖTj�J����dG��X �R� 	`�+p����KIɦ��P*�m\�T��z+T�⥉8!=S:�n"��m\頺��k"�vB�*UO�zJ;�R�4���Vϔz��<!ߣ�Ki�V��R��Vo��[�8�/�x)�Ki�V���n����n��}UJ�R��<G�UI���u�.*uQ9ή�Ee7VI��qv%%*˫ʩt%�)���Au��UYqU������Te-�D���R����v�����e��*�O�x&��l���T��)�O9���?eU)�&r�<K�3��Ȯ-EP9��DB�*k�JT����URq�m�*ۥ�v����%Q��)�O�U����c�ʮ����7��)�M�U6B��>�����45�ظ�Ԕ���W�FM�"�0���]��9���d��8%�)K�ʒ��$�$;e�SY�T�����9e�S�s��r%�)��b��ةlq*O��T*����T<e�S��TZ�������l*OY�Tr�\��T�3��L��)O-��r-���c��б���?%�)���b�	���&���J7T��rP]�U6B��Oe�Si��ʦr]	����ũ4H�A*+�*ܵ�3��l^*gĕ���E%%*)QY�4��������楲y�4H���CZ�TJ�R*�R�4H�A*�ҕ��,v*uQ��4���+��G%8��E�U�� �%Q��� �i"W�CZp4���zy� ��,�*YRɒJ�T��+�R)�J�TJ�R*M�|�o�vP�xi"?�ې���L�g*ۥ�iy崼rZ^)�J�TJ�R*�R�l�*R�AUvP���J�T�K�UR%%*�ٕURq�4H�.*K�Jp4��w�
�J]TR��]��;M7TN�s�&��ӓ�R���c�U��O%*�J$T�8�H�DBe�S��J$T"�:>X�l*EP)�&r�4_��z*��&�B��TR�����E儻�8!)Q��4��w�J�&��n>;���	M�	�h��n�DB%*EP9ήAyU}���&�}i���Je�RI�J7T�������J�S(�Je�R�����L��ӝ��)�͕��&��n+�͕֧AW�y�Ae�R��J$T��Dw�"��?��)aO	{J�3���]��)�OټT�,�5K%*�P9-�,c*�P�J7T�1�����W����Je�R�ʶ���^�m���,�3���R*�R��;�R��J�T*�RټT6/�#�ʚ��8�ĩ$N�g*��S�J�T��8��K%q*=�D~�w�SY�T��R=���L�g*�RY�T	,YR٩TJ��<���%��He5�D���%V�TJ��K�T��+Ri�ʚ��f��Y*R٩4�Ku׶|���J�*�PY�T����qX�T�%���JpT� ��G����8���CZpT���-�lK��O�QnRكT� �=HyB�!�J�T������E�.juQ[T�R����-*j�Q[T�6	M����E� k�P�Z7Ժ��oh�?>�sdM��⭶G��v�]k��&���GmQk��r�� ��5H�AjRk�Z�����ǆ�������>����r*];�n"V�j�ҵnhi\k��ڠV����E�T�V����jk��ڠv];o�eIm�P˒Z�4��Х� ��-�8��%����ڠvP]+�Z�Զ��,�eI-KjR[��V����p�v���ڠV*�C�Z��6	�x��K턻��8����UO�zj��Z��v��E��jmT;��Q��j���V��8�ĩ-*j�S��z���3�EE-qj�SK�Z�ԋ������D�B��<G�ڨ�F���k��D^Bo�/��h���X�����h�@k"��w��m�a|��j5V��Zz�:�VP�����ע�v�^���ҫv�^[��j��^�ΪuV��j�M���M�F���D�&���l��Q�佶J��j�W��Z��b��q���5[�T�&��Y�Ϊ���cy����zj5V��&��nw��Zzբ��ةuV-���������Y��Oq����ExPc��QmoT��N�k��D�or���Dw�꩝�ת��8M�o���ꩭlj+��~���i"O�/��V=��UO�Tw�6j"���b��\����ݮ��Y�]Om�S��4�h�S���~��j��ڑ}-�j�UK�Zz�ҫ�Y�ΪuVmeSK�Zz�ҫ�^�]Oy�>~���v=�]O�����^m�S��Z��2���i"W�@��v=��k"�v�q�]Om�S��Z��b�{�ث�]�욈E���F�������F�ث���;�ث�^m�T;��%a��j��M�"�O��Z%֒�������jW˸�9x��Vv���e\m#T+�Z�5���J�m#T����v�^;@��zj�W[�������-vj�$��_m�SK�Z֒���u�Ub��j��k"���ث5[me�D�C~hʮ��n>�V;-�5[y,��j�Vc����W�h��^u���8�Vc��M-�j[�Z��j��^����W��U���Zg�r��F�]O��jmT;\��Qm�S˥کt-�j�Tk������D_�T�ڨ�F�6�T�r��K���ڒ��$��zjU;ᮭj��qv-�jK�Zg�6B�Ϊ�zjU+����v]��4��� �j��&��(�j�UK�Zz�ҫ�j"���'l�j'ܵ%Q��j�V��2��J���7���k��Q��j��$�%a-�j��&����^�T����v#;��5[-�jg׵f�5[��j��D|��/Ď�k�&���?���Sm�T3�.��^F��%��F~���ݵ/��Xe�	���y���k_�~�^�"~_&�}'����Z�"���ޞ�wo�����+ً<����<��;�����G���8����e�E���>�"/��+�D�_�_�������&�"O����E������\��k�D��^�?�}��'�M����B½������~�S�D�:�q/�����^亼�@�&�}Sx��򞃪{������5^/���a�E޻	^�E^U�&�w���c"o0����K����"�����E��;�E.��KƋ<���ʋ<�w&�ދ��ކ�{���6D�؋<��ɋ<�w&�ދ8<�E��"~h���ËX*��E�]K�׋8G��Dn���r���"/�	�"�e>ߋ<����"�����E^{7�E~��ׇy��_^�?t�a�^��i��.7T�E^w-��%6��
�"���0�
`�q�To������û;�_/�"�&�iE׋\�{��"W�2��^�����{�?Z7�k"`L�{���G��E��z���i��z�M]֋8��E\{�&�i�z����h��k�z�K�1�W/r��G�Ջ\����"?�g��E~�o��{����.f�E.�-��z���K,W/����"/����"�e�ދ<���h�"O��Ob/r]>�`\/���k'@�E�C�֋����yxw-f�E˗SJ�^��}"ø^�Rݢ ���^M�S��z/�ݏ�G�q�!�^�/��
A�"?��EX/�����M���E��{q��{��gz���j"sx�y,�1H/��z��v2��E�C_����G�U/��q}4��&r�0��E^U����^��'�s�1�z���c���y%|�^����z���3�"O�7Ql�D>���"��ӊ	w/b����T��^�'���7Q&ܽ�J72��EލL��D>�h�z�'��`T/r]�:�G&Zy��T�E.uY/�)��^�	y�@c�ȫ�}���yq|��.�E�8���FN72@�E˥��
�z�'���"�0[/��X/b ���r��g5�o�����"��M�>���� �yx�6�E�]�Ջ����AU/���~,���yxw-��E���m*�^�|���^�|��E�˛S�&�>�z��� �z���v�q��O���z?G4֋8<#�&�{m{S@cM�.�"��ӝ��k��z��p�#�^�|"S��"��۝"��܏p��߶���"?��z���@���nZ�&r�0y�E��_u�Q/�]�G]֋~O�K}L�{��ir�O.�Ѡ��ߋ�1��E�g"����W����Y}
�OA���5[��F}�q��c�����z�W�-:���J�D���=�S=}��O��Q�5�̏���؏EX/�z���dIyB�ڏ�|/��<��ϝ�.��ȶ}��Op4Gp�I�>)�'�DB�H�g�E~"ﾟnh��E�)�z���e"�D<E?ڸ^�'�E�E���}R��\ߑ?��G�׋���m��G�׋�8���@]���>)�G�׋�D�&�����y,o
����{�P}�}�G�׋8��裳�E�'���c���<��Zz�^��Z�'G'�=z"?ѽ����'8�h�z�K��A�[�Ku�j�>�G��D�Z�ѧ���?m޶?�^�Ǳ�	����>)�G]�D>�)�z��w�1]�E�MU��e"����4U��s���E�˝FyՋ\���{�G�Ջ�Dw�����E~�OdN�9ܵa��E��i�z��ލnQ��^�Ǳ���Z�ӧz�TO}V/����B}z����/r]|m�����ɐ�y%���Q^��B}�Y���3}z�O��Q%�"��O�M��J�E���L�q�eI��^ď��{/��Vz���|/r�4��D�/�4U��+�~���E��[�)~/�XnQ*�&r��A5�V��x�V�O��	�>����qB���)~/��h�&��>eI�R�0�%}�K��k/^���aH�ԋ<!�6UR/�ݵB�O�1$�E��]����c��(����r��v��Cs?��>Qէ����"ﻯ���Y}:��v��z�^�'R%�"�%Q/�z17�E~��X��"O���f�]�E��7z�^��}n3p�E.�;���Sv}tP��O��.���T8�7��@����>��D.����SvM��)�g�"��}B��i���MA���>j�^�"�K3_�ᩥz�-����z��+��UP}�|WU��)�>��Ǭ����xi"�����DM�O��i�>��^�R�%�]�E��h��Goԋ<��8}�O��Q%�"��[��ZY�'K����"_>��K�R�S*}�K���x飃j"�\�g��K�T/r]>��K�R/��X����a�z�TO#�^�i�|�K}r��Z��z����OA5��𞣳�T�\�K}r�O����>�ӧz�$N���c"���D�&�W��������E~��!!�GyՋ����+���z���=����zj�^�	yϡ��E�8(�z�������R�SyS�K}r��\�۽}-���E�]۾���r��^�	�T��^�"|Hk�>m��D��T�UR/��%�*�eo��3-=��3-���w�K���KK��8�"?�m��zZv=-f����u����i��K�"�ʣ|	��jY��Q˒��<�yx��.{���j1��E^{��KT��z�"��c�㦰�X�v�e�ԲJjɸ�fki�&����kɸ��kɸ&�7�{β�j�A����"�e-ղ�j	��_�"l�Z����Z�K-IزJjY%�$aK�d\KƵd\K����"���}ɸ��kɸ��Q˒���Z;-��Rc-���Ǘ�%�Z�%�Z�%�Z�ŀ�y	y�_�^|���;���s�묖�j�⴬lZLP|KUcM�'���k1Aq"_�o
ҫ����k��Z
�e��b���8�Ku?ʥ�_��}�Zƴ�Q���/��X�����yx�$�l^ZB�%�Z�|�K�1Ǭ�q�p+0��E,5�%�F-f������RP-��R=-�Ӓ8-����iI���iI���hI��eL�2�e��� -uѲyi	���KKp�Gy�>a�=�TZJ�%KZ�3-���,i1S�E˷�p[ɒc�^�'ʒ�i"N�z�W�� ��z轈�>t,cZ�1-���3��sH⴬lZ�,-��R*-��bދ\�;�N��<GM��e��R-���Ot�	���K��%KZ��%KZ��eeӲ�iYٴ�L�~�e?ӲSi�s�^��-PZz��8m��D�Kϴ��"?�'��iY���K�9x/�X>��J��x/�X>GKp��EK]�l^��+�� -�޽�O�S��lqZ��AZ��AZ�u�V��{�?Z��v=-YҒ%-�-f�Ų�ii��iY��dI�qv/r>X5H�F�%KZL�{������PKp��D˒��.Zꢥ.Z��%�Y�%�YZ��<mw�]O��`U-Eв�i"/�V��b�݋�D��v=�WQ�w��~�����%%�ȥ�E�z���^]�DB����-����&r[������ʦe?Ӳ�ii�&�����K�楕>E�J�qv��YZv*-=Ӳfi陖5KKϴ�Y��O�)�gZ6/-����iYƴ�JK���J�2��\�ٚ�e���3-k���i1��E�C��M�-��L����ii���JK��dI�iy/�zټ��JK���JK��dIK��4HKp�GKp�GKp�G��w/��0�E~��т����� V6-+��,iɒ��KK]����"��v�yiټ�4HKp��D�	w/b�R����ک��EK]��DK$�A�Au/r�>~���HK�3����\���P$��TZ���ZL�{�Ku٩�7���)j��R-���^�R�0�{���+�nh���Hh٩�DBa�R��N��S)�T
�Q�©t�A
�B��pv]ȒB���p�](���/���B��P*�R)�J�T
�R(�B�v=�]Oa�SH�B�z���)�L!^
�RȒ®��%�,�5�znC�"����s;zN�Y�+|4��<��F�P��Pa#T�B��?�"(.����O�������Na�S(�B��8�-N����'�y��D�+,c
˘�2�����'�g
EP(��ʦp�[���㜑�r��B7����7e�"��;�3�BJ����)�Da�SX���P��N!8
�Q�B7N�����ra�SX��p�\��b�� �]Oa�S(�B�ΛYRȒB���;����c���8��)�
���t�z
GЅ�P���F�S�B.r��K�\*��
��BAVI�*AVI�URaoT(�©t��
�{s3���
k�Bg:��Y��*��
��©�m�<�7���
�B�N��yx_ӭ�
��&��:?�C�5�WշIXX%b�{�f+4[��
��D^	��_�C����p*4[a�Th��*��l�f+��
{��zaoTH�BgVI��j~/�^��t�B����j"�Y��R��Tᘽp�^8fo���p#�z�^�p,l�
-YXK5�����MUa-U�B�b�PvM�ܢʮPv��+d\��
���
]��v�k�ʮpZ^X^5�?�m��D,U867r?��J,Tb!�
˫��\��]%6������¦�������򪰼j"O�'��,�ea�U(�&r~�w�_(�B^�^��,�d�%;���~��X��B%���p*��7��ˍl-U�B����W�T�FM�|H[%Ne�D��w�|	�W��B��F��QaoT���!�a�T8$0�d!�X�����
g��$,$a!	�W�N�XX%VI�p,N���Bq򲐗��,�c����*�
;��!���H�	]Z��B���pn`870g!/yYh�BKa��,�d�%���EX!/�X��{��U��
�W�g�Y��+�^��
eWX^���W�B�b���j">�|�U��Wa�U��B����*,�
e�D\	e�D�/�����*�]a�T(��v��q��+�����<�C��@+,�
�Vh�B���h�3�B����Jj"Oۍ,�
�UH�®���)�����B�2�h��j"�ꄻ��)4[�ٚ������)�z��1g�S8/�]aS8�.�g
5�D��0+�B��Nkw��+�]���u���>2�
�W8y/�^!�
�W��&r�>Em�
K�B�b�{m��v���m���m��v�ޖ�mIؖ�mIض�j;yoǶJl�ĶJl�ĶJl�ĶJl;�o"��k��M�Ry-�vcmyٖ�mI�Vvme�Vvme׶�j;�o뿶�k"��7��V\mIض�j"?�7�-��6Um�׶�j[K�%���b�m��m���R�Q�[%�m��*�-	�	ܒ��<�7�ضjǶpl;$pkɶs�pl���c[8��c[8�m�ږDm���P�F�-/�ȥ��c[8��c��c�&�kUb�©-�±-۶Km��v"�v"�V�m��D�]k��{mK��%Qے���������������ڶKmg�m���k;�o;�o��&��xX>ʅc[8��c�>����<��$lK¶C�$l"?ѧ��>!��em�ضkǶJl+���k[��%8���-�|H[���_[���^����-���w��v���m���k����k+��Z�����-���lm��D�-nQe�Vvm�ne�Vvmזqm5�D.�����-����^���Wz�uVۺ�-��ҫ����G��m{��@k�/͚�m��vH��qm�D,�+a�D�����ݵvvm;��$l"�Q%6���U�mIؖ�mIؖ�M�"�ے�-	��E���ے�-	ے�-	�b��<���­�ڶ�m[¶�k[�-�*�m��vx�v,�֒m���m�׶�k���]۱�y%�u�&�����Z��%�B��%�±���F�֋m�Ŷ�b[8��c���l�����|�[/�Eh[��g[q�g[^�-!ۖ�m��֒m���m�׶qlK¶$lK¶�c[�%ayB��_�Ub�z�-�*��ێ8�*����m��֒m�öplǶ]b�.�-�±-�±�ksql	�N*��mK�֒M���i���8�֋m�v�ᶄl�Ҷ�d[�6�4�ޖ�m��D.�o庴m�ٶ�l�Ҷ�e[��m/۶�m�˶zm��&�c���	Ͷ�mڶ�m�q�m�j��nb�ٶ�l�^�g�و����K�"�-B�"��\�_Dhq����K��Y�V�m�ڶ/mڶ�mڶ3��jy��MlU�J�-{�����{��m%�V�m��&��O88r;%r[��%t�)��V����Dh�b��o[Ƕ�^�Β�Β��c��!��r����ڻ�������xɭ��Β�����n��n;qr;Kr;Kr;8r[ڶ-mۖ�m��V������ֱm�޶�m���m[ڷ�}[ڷ�q�j�mCۖ�m�?nڶul�:����j��\�w��vp� nK۶&p � p[ڶ�%�˻��$�Lp���m{۶�m�޶�pK��p�'�B��#9ܒ�-9ܒ�ms�D�˹�[�8���f��vz��=n��V4nGUnE�V4N�9zKsz嶾n���q;�r�{����.o|N����m{�%wے��ǜ�E�%�ܶ�m��v��Vmn��hN���'����m��_n�vn=�vh�vB�no|��m!�Vmn�}n!�v��v�綵o�6�s<�Ds��:��#�<��#�<��#�<6�)�/��
�(���(�|�8��('r��s��w�޻��D^��:�#�:�#�:�������xG�x��޻c���Ƿ�#�<R�c���=�q{��H!��8��#�:�8��&��zǩ�ǩ�Ǧ�c���P��L��q��i�8hs"�����*��7���(-��}GVyd�GVy4�GCy>���c�q�U+��}Ǌ�#�<��#�<��c��QGu�QG��9�Ͻ-r��u��>��:�X�wԑg�k�;�#�<�ɣ�<�-j�ݑB)��؎wԑGyԑGyԑG�x�y�;��#_<��#_<��#_<�ŉ<m�������8�ءw��G
y��G
yl�;V�M�'�-�h('��p4���c��q
�_����QZ����D��|g�=�D,B�y��G�y�㛈+��<����Qm+����9�}G�yT��־�\��![���}G�y��n�ckߑ{N�'��� =v�Q�D^h������u�n�#0��uy/��hNO�������cO��{��\�~�Xx$�y�������D~��/ꑡꑡ'��q�q��q�둎g�5�s�I'r��`�!<����أ9=��c��q(�Q�5鑎�葎���d�u�i�G'z�Gz�yx7��8:�8'�X8���U�5�qN�M�L���_W�G`z��G:zt�����=v��s�HG�t��9xt�G'zC;����)�D�(�(@��� �N��}yЉ�豙��LxԤG:z�<jң&=����ڣ&=��cu�D�C��Ow5�D�����;�Sn�#m�#m�2�XixĪG�z4�Gs:�'�}�J�#V=���qX����+�9=�ӣ9=����p"?�/�#0=V5鑎����
���98��+O���u?�=�D�H4'�ݢBΉ�D����XCx���6�c��M�9�m��z��t"���~�o
:ѣ=�=��#=:щX�e�G'zt�Gz�ǉ�s#�}n�=����_x��G�9�K�����û�U�G�y$�G�y���J��H�#�<Jˣ�<�c�Dˇ���#�e��1�G�x�!<"�c��9��Q4��Q!G���c���G�x,��E�LS4��Q!�Q!�����&x$�Grx$�����B<*�#9<2�#<�����*
 ��o"���9��Q�M�"|̕�9M� ��M��M��M�q���� �߱��H��e���#�;r���;ڻ���#�;�=ڻ#�;B���;�U�%ܑ��۱���Lx�qGw4ny,�D�!<�c��M�8M�HՎT�HՎ�W�v�j�6�k���JծuW�v�kW�vm ���]+��z�JծM{W�v�jW�vuiW�vuiW�v�zui���8���]��D^/��ե]G�^���T�JծS[�z�:i�*ή�V��{Wq6��b#_�U�]yٵ|o�?��	)ή�l"���l">�־+B�"�+B�"�k��ե]��U�]��U�]��U�]��^���.��Ү.���&r�ZO�"��8`���wEh�n�kkߵ|��ˮ��jɮ�z�I�WK6���]+/��%�����Չ</��I��Z�+�v�]-�Ւ]-��]k����
Ǯp�Į�V�zWKv�;MKv-̻�U�����C��]]�եM��O<W�v�[T�v�jW�v�jW�v�jW�vui�y���W^v�eyB��_�ٵ��*ή���ˮE~W^v�z�dW8v�c�"��%�Z��%���kE�{]��Uv]e׵��Z�w�_W�u�zZW�uZ׊�kE�D��w�D�����k"�C�u5[�����nd��u�D�8|�^]���Y]�յ�� xEUWTuEU�����k)��^]K���:�����몱�=�W�u�	�����ʮk��ut�`�꿮m�W�u�^W�u�^W�u�������kO�Uv]eוq]��^e�D~��e�u(�u�'p"ወpl"��@%v-����p�Į�d�$l"���&x�_W�u�_����ĮJ�����d���]�J�Į�d���꿮Ձ�x��M��O迮=�W�u�_�ɴמ����uy��]�ص`�j�&r]ކ�cW%v��*���+�±��D�`�cW8v���O��x7Q�]yٕ�]-�U�]��U�]Iص��:��Zi8���;���!/�Z����+/��k��ub���Ү.��Ү]������Τ^��Ex��M����uyS�]��^�
��ZV8����½vN����ǽ6^A�U�]k��Ю�Ю��&xEh���W�vEhW^v�dWKv�dW8vUbWv%as����+	���ku�U�]��$�Z
8���_86�PKv�dW%vi{%a׺�k�ߵ��j�&������:�*�&r]�Z{'r]>�-�R��K���k�p"���.h���k)�ո]��^{��|��W�v�{����ڽJ���8�-���O��Pnw����w�u׺�+��������^ �3z�����uWw��佶��r�K�E~WUwUuWBw�r��׊�kEߵ��Z�w�v���mg�^[��h���E~W�7�����]���]��n�j����]����h7��r#+�%wq���]{�%wWUwUuג������k��U�]����]�_���t��kݕ�]9ޕ�]�	_��h�:N����h���h��h7���@�wu|�F�k1ݵ������J��hϩ���K_:(8�})�K��Ү�tPpj�F�t*p�S&�� �%w��t�o*S9�����.ń)&L1a�{7���w�T�]u)L�`ZL����� 0�})�Ki�D.�����.-���E�����T��ui}]*S����8�̧�/�ћ���.��2��	�L0?�R&�2���/u|���z��K��B/z��K�]Z�r��&.zi'\��Қ���M���v�/���M�Uu�;�7��K�`~nw��D^���u)9Lg��
1%��/���{��G���O��޻��.��i�]�{��ޥ��S��Vᥳ�Sј�Ŵ�.��i�]Z_�N�Mb��I��$�t�oZ����T!��0%�i^
 S�j�T���`1]ZL�ӥL05�i�\�S&�2���.e�y%|n;�7ۛ����&0�) L`�7�N��<��m�`*S9���T�L0��K��I�)L�`�'r�>��) L�RڗҾ��M�R���ֱ�&0������N�����NM`Z����r0����5]9���T���S�
�T�/�xi�ZJ�RB�6��MhiZ���r��Х�.������suSB�z��˥^.�����Х�.%t�ݢ��Ek��ݴh-Uui�ZJ��V��nQ��Rh����h-�v��K%\
�ҹ��qK�[Z��N�Mk�Ҏ����-���֞M�'�`��,5ni�Y��R����M�[j�R��<�;7m)hK��&�}"���--G��û�m��Ը�z-�k�ݴ/-5ni_Z
�RЖ���	-�;����R����-5ni9Zj�R��Ը�z-�k�$�T��z-�䛂����}Ӣ��-�ei�Y��҉��xܴ�,-4K��N��?t��4-Yj�RK�Z��/-�ci�Y��R앎������MT�����������M�%t+XB�6���b��t�lj�R8�±T��]bi�X
�R8������$,%ai�XZ/�v��]b��Ԓ�Jl"W����J,�_i�X�8�N�MeW:�5�])�JK�Rٕʮt�k*��^��<�����t�k*�Rƕ��f+5[�}h�S[ӎ��q��+mBKWʸ�r��q�MhiZʸR��֞��\Sٕʮt�k:�u"��*s���,�8K5V��R��֞e�E�wL�Vj�R�5���S������j��J�VZ������k"OȽm9ZZ��2��--GK���r��-�=K�W��҉���J��D~��X%a�s�h-������h-%a��J��R���CNS%�*�T�e�7d�XJ�R�ʮ�q�ul��JWʸR�5�B��w{��ҶTv��m���{�#GS�����$,�vKG��J�$a%�*W	����l�@��q+�V	�J�U��~ڥ�*Ǘ�f�4[%�*�VY�6��O�4[������ny	�����]e\��J�Ub�r
i��>1��������k"��ޞ�ճ�˚�{�5qeM\��ʚ��&��UZ&-������`�Ғ����+-Y9���^eM\�J�UN!-���p%+��D��;����d�%+�XY�V*��<����`"/�J^V�-yYi�JKV±R��J�,�+�X�&�X��]��p���J�Uʮ�q�f�4[es\�Wj�Rc��j�[s���(�*��JzU�ĕ5q����ֶ�U���,�+�UY W��M�"|H��6��p�Z�VV���ne�[)�ʑ�%�*eW)��a�%�*狖���]��*eWɸJ�U���l��>K�U�h�@�Z��; ���YV���n��*5�D�g����Yj�Rc��7K�U6��m%�*�VY�V��rgɸ�����l�#4�:�
w�ΪDUe�ZٽVҫ��D7�@�tV��*�UY�Vҫr�eI�ʆ����lh+�e�ule[Y�Vֱ�ul%����h[�&���o���Ek�+��J%V��Ek%+�XٽVv��p��ce��D���-YٽVZ����$��K+�WٗVb��q�}ie_Z9U��K+�W���
�����=+k��ڳ{��ge�Y9	�Tb%	+�WY{V��r�eI�&�-G+��J%V*�R���2˾������=+k�JV�����ge�Y��J%V����$au|�ۄV6��p��c%+��JKVV��j�8+yY���q�e�Z��J�V������e%/+�q���Y"����g�8+���V�����Y��ҥ�Ek%B+Z٪V��ҥ�.�ge9�D����i�e_Z9 �4ne��Dޛ�Ek%�+q\������+�ʆ�����c+�]��V-K�JhWB�ڕЮ�vei[9���q+��N�R}�~��� I�ʚ�R�M�"�3�	W�*-�`��渉\�/[�=-}a�˹�������Ąe1]Y97�N�Ǳ8!�aI�������ҿvZ9Wb���p"W�ILXb<�����,�+}a�K_X�²�n"���b������+�b	K�XNG-�b	K�X�ɕ�қ��re�\i�ʹ�r��וto�~��_n"��ՉX����e]�K�8���/"�Ĳ_���e�\	���U,+�ʩ���5iK�Xr-��ʮ����D���rlY_W"ǲ��t�eW]�UWRȒB��t��{,�cY9WVΕȱD�%r,Gǖ�t�eW�D.�[��ue}]Y_WRȲѮt��{,�c��޻�Ѯ�Z���=�|���e�]�hW6ڕ�v�h����� _,�b�K�X������	E������'�+�c��F��=��ty,�"ǲ��D�%_�ȥzSho
��M�O������.� ��R4���m�k��Z�غǶ����k�c�U�R��=�]u-rl�c�'򴹛L�9�%��k�c;�i�ӵ�t�{���{B|�h)dK![��ίm�b�h׊ƶѮ�k��Z���Ŗ/�V���y,�Bl��Z��*Ė��%�-9l��Z��ӵ0���-Ll�ж
��L���&��vy��Zab�ۙ��4�&��v�Ul��D.l^�[��"ǉ\=�m�^�[����M�R��X�׊ƶ
o�'���',�k��D^/o
�vbn�U�ӵs[�غǶ��u���ܶr�u�m�\;W�u�-rl�c��Y�m]�B�R��=N��?���"�9�ȱ��k�c�B�R�v�mK![��"�9��s��V4��j[���Ķrn"��C�1���p��[���m��Z��"��*�erm�\�2��&���mM\[�8���t�渶9���-9l�¶Caۚ��&�U��Blk�ښ�����4�b�׊ƶ&��-_l�b'r��4�'�ݏ���*�0���mM\���*�
�-�kǽ�
��[T_����N���Y�]uq7&�0���m}]�����]u-9l'���
�6����m}][_�ZŶ�����Ul��Z����vl��b��*N��}C�/�|q"?���]u�{l�c+[�8�����hl{�Z�8����!rl�c�[�؊ƶ
�E�-rl�c[�7��ض�m�k��Z����=��E�-rl�c[��"Ƕ
������k[��Z��*�Ux-9����7ab[��Nmmab�[�����������޵����޵�p"ወ
�U�m�D���"ba^k[rؒö��U��l�v�k;۵勭Bl�aK'���`�7��F�8�W�{�0�%�-9l�aKۡ�-9l�a��גÉ�~aQ!�
�%�m�_�[���<���`;`�ń-&lgζ��ńma�	[L����	�L��!lM` [ �N�m'Ӷ�-l�`;����-lM`�L�6�r��_�b¶��ń-&���{�v��G_8�ڻ��j[&�:�����q,��;� ��?Y8��5��dږ	�e��ږ	�L�m&���� &l1a+[9�2�v2m[|��-��/lGڶ�K"�BlbK[r�N�m}�D�C�����Bl}a[|ض��j[_�b��]��l���*�l��D�8�*"l�`;Ҷ�������ͧ�k9^��Z��r�ڵ5�ma[C�r������lU]�&�B�ڵf����X�5�-ڛ�u�Eu|��k9^��Z�׶	�m�-�k�]���yھ�k�Z{�Μm9^��Z��r���ch[���m;[��
��޵�m�`;M��&�v���x-�k9^[C���h�E{m3a;�v"��s���H�����ct����>�m�~� /r����_�'�>�_�	����������E�>�_�~oC/r]��yq~�L�{�z���}-x�W����"�W�7�����������<��?4N����"?����"?��>�"���1�������7��;�{�y�K�����u����E.��n�"�{�y����y����u11�E,���/r�Sx���}�y���f�B|����
r8����{��/򄼛 '�}�y���_�"B��>/r�s��/r�/5/rެ��"����D�:0���b��ջ�i9|��˽�	|���F�q�cX�8�r�-��~/�2s�E�6&p"w��E���Dn>���<!�0�yB>ʑ�/��~�����q"7]�/��|N��C��c�Z@��\����_�|nc_��ݵ��y%�| ����5���E�>|���p"��̜}��(rp"��`�q�Í�/|��poC_�|�B_�"���ĉ|�҅�"��۝�ĉ��(��z�|��1�E��v��_�'�k��������<!�(̈́/�� �q����q,.!r�E�6r�E.��/L�E�˽�	|��roc_ą��p"�(&p"7��E��{h��y�E��;��"?�mE����8~GF��ջ�@{/r~��s�E����Ɗ�{��p?b�������".�E��E�#=�/�����V��zw��E����{�K��
�{��Ч(�d_�|>R��?�9���}"�xR��"��/�n"�x� �"Oț=�/r>��|����{���}�R�������"�����^亼���"��k�_亼��&����^�'��^�'��^�oSn'����������"���B�E����������^�"� _�'�-���y%|��s�E^	��_o|���o|�	���.Gu��<�7+�ߋ�8޿�	|�W�;��_�'z���E^o���T���O���E,�7�9}�a��8G݋�D�#8�E�-��u���"����^��V4��ջ�z/�����E�C��)��^����<��E^/_ t���"��p�D�����"���E�	�"~i�{�gP��<�[��/�X>Xao/r]nd$܋�^nQ$܋\�V����c�E�{��>ao/��2O�݋<G�(%w/r�>i�{���w�r?��^�9�wrT�D�G�݋\���pz�^�|���^ı�w/��ؾZc�^ą�޽�sڽ�Ex`���Do
����-�A���@�ދ\�w ߋ\�|hߋ\�w�ދ�D����|��޽��}U�"���n�۴�M��U�"O��v{S�˽�s�����r/�=�O/�ю����J���_��(�{���S�}�O�6��ɧ8���{��bw|�Ľȫʆ���"�O�O��Q9�"�s��M�'����k�z�S�}R���/��<�?�٧8�g��죅�E�����_���{}b�O���B�"VO݋8!�ا���{�K�Y�I�>��^�Ǳ��}±�������c�v���c���_n"���q/r�nwj�&r��Zj�^�o���p/r<?߾���j�	�>��N�S���E~"�Ǐ���	�>&澈���">Qq6��KȨ��ˤK�ti�.�ӥ}������.^�?���$����m4ڽ�Ot�K�>J�^���q�.�ӥ}�����y��Dhy��+٧K�Dh���S�}���!�/r�|��Dh�t/��GO��|��h�"��C����>��'{�do��m"��p��t轈+��߉���O����>�ڧ^��j�}_ď�I�/������O�AxSP�}4�M������{�>����yx��1��E^	o
��M�k%w�ki�{��p�2D�E,b��v���}"����yx�����/�}֊�>�辈-*B��{��r[m_���"�ꃕ��/r��Z��>Z�^�|����E�ͧq���{A�'h�m�å��e��\��G��^���|>m�T��}�M�wQ-٧%��d�j_�"|_Ւ}Z����|��}L�}���q"��(Z{����S�I�>Iا���^���{}b�O����>�^�i�
����_����}b�O����>��Giۋ\�VI�'	�$a�$쓄}ʮO��i�>��'��
�"��|�R��"�V��I�>��D��o�ҫOz���>Z�^�R��ȥ>��G�ڋ�D�&:�OA�1�u"�;�g/���ڨ���y%|�ʥ>��Gڋ\����Tq�r��ڳqx��^�	ф��?�9҄�"�2�e/r�>��:��OA�1��E��/�����c��PT���>Q�'���8{����j"?�-J{ً�D�j�Oz�I�>��G/ً�	�DU}��OT��8�"���^}ҫ�.��.����#�J_��i{��諵���Y}:�O.�Q�"W�U}&��]Kq�Dn>է���Ry,�⧠��R�\�cr��D�U���Q��^�E.�=$���P��B}��O����>��Ǵ��ڨO�i�>�ӧz�$N�a���L�j7�c/��K�>�ҧT�(!{��ޯ���z��|dʒ>Y�'K�dI�a/�c���G��^�'����δ�y�nw���s����/��uPB�"��\�K}����yx��ڨ������'�=�e��b&��D�1�/���,5ֲ�lY/��[֋-��b&�<G�/ǖ�kY/��[b�e�ز^lY/��[����Z���,�b��<�KƵ�%[2�%�Z��������n�,![ʮe��{-�����&�z�eq��M�'�ֱ,[�����Jl�ĖJl���J_�U�-��R�-��R�-IزKl"����bKK6���f�%��E���e��%/[�eU�R�-���Q_��y�Y�%/[�����ކl��O��g1��E^^}��I��r�"�F��Dh���Ŭ���������������zy�Z�gK8�$aK���U�"W﮵�l��&��ǖgKK��8[±e��Ғ-kϖ�lل����"/!_��.m�Җ.m�˖�l�˖�gyB��(�&r]n��ޖ�-k��Q_��r�+Ζ�l	ǖpl"h|aYZ�%	[�P}�(	[LZ}'$	���{S��P[V��v��q�r��%[Z��%[Z�eڲ	m�˖�hKq��dKK��dK%�Tb��/��n���ψ�yB�m[Ֆ�l1��Eޯ"���K[v�-��b�닼8�`��]_�"�v���oC�-	�<��^ޙ�[v�-;ᖝp�N�e'�R�-k�5q˚�eM�R�-9ޒ�-FǾ�uy��n���ho���5qK���&�"�-�2���[�}�?_W,�[:�%�[�����z�9��n"�[�-���-�ޒ�-��Ca_�	�FǾ�Exϱ�nY_���F��	\����Do0��M�'�h��"��0�E\/�떘p)�Lp�#Z_����_�����rpY �d�K8��蛂 p1|�E.���<��*\2�%\2�%\��e'��.� .��&p����oI���o����o���q[�c}W���E���ҶŤ�q�j�ei�D~��]��^[v�-�ז�oY�6�����oY�����"�CZ&�d�K&��^[v�-���.[Ֆ p٪6��r��Ą�V�%&\b�%\2�%\2�%\L}�'��.ږ�p1i�E�ˆ��/\b¥\�v�	.���	.�ݖ�nq	���p�	��n�j�%9����Nn��&.a�&N�"�)���p�.� �,�K���[��ň���M���渥U\Z�esܒ/N�	��U\Zŉ�8�ǛBzS�*.���ȋ��P4.���q˚�eM�b`�8!��LnI!�rI!�r�B7���:rY9�t�yx72sO'�_�8����mM�D��܏�ȉ�9�Z����T��-tKV�4�KC9���~���l׉��U���Ki���KC�4��2����q�v���]V�d�KV�d�KV9���>a��b���D�{���[�ˉ�D_l�[6�M�Ǳ�8��/��qK����[�v��?3�1�]_䯉�=��c.=�b��\�����#�\�h}��ro&�`r�/���"/����_C�ԑK��P4��1���t԰9.���P!�&0���;�&r�쎉~�k�����-d��	M`���*�`(C&�*�B92��	�SHC&2��.d�����Nıl��`89t"��_h�B{����.,m�]�Bh����.�v!��¡�aC[��BU휈_9�]8�3$t!���c�kUu!�	]��&�y��3A�N��x��]894��k�B����CC��ą5q�|�p�hX&j��L.�! ` �ʹ�r.4��	M`X92��\��`�C�� ��/��`��B���P�B/za'\�	�����)��B�����i{r�i��B�7�K��z"/�7+���b�P�L0��`��b���.l��`(C9V΅�s!&�`8V5Ąa�\�	�ʹ���0d�a�\h'�J�B��p`j(�ʹP���r! ` '��F��X9����&0���-ta]8V5,��`�C�Ҿ�h/l��]�B���r.Tu��U]�UvՅ]u���\��B/6څ�.$ta�]��B/z��˅^.l�	]H�f;zq�X�B�P�M��'�-̛��{SPՅ�]CB�ㅪnn9^	7�^.�ra�]�����и�zm"������u�^�B��c�Z���F�ХM�"�;�*�P��z-���ׅ�u!h瞆�-��[��B�NG����y���B⸰Co"���¼��M�"|�J�BVᅽw!U�ZX_�ׅ�-ma}]h�B����.�k�^g���-l�g���JC��ޅ�-,��[��B������Uxa^X�7��������G��v�pVi��BB��Ѕ�.l�U]��BU����k�K�6����&���;�4zak_��B�r��ㅣP�Q�!��^(�B��B��D^hoir����.�v�t԰�/�w!������r���M�'zg��3TChv���~!��]h�B{NZ�]��BU⸰0�ra`H�BB��0�q!���O�`)`X
6 ��.�v���� ���p"�Y��M�"�O8�5z���^(�&r����B��Bo"oa(�B�ڻ�ޅ�n�?�M{6N�'�9^XV
�pl(��f�p�k�L8�'䋈���P���&0l9�`��B���ptl��B����h/,>��i����_H�B�:�p�lثΜ`ث�*�&0�a�bhC����&04��.�`�C&��pXm8�6�h1a8�6����`X��;��0lr��s��Gr�Ð��kC�*İ2V*İ2l�abC�*ĉ\�oV��&�01$�!9�$�:ɉ\�wL'��qâȰ(2l�Ec(C��ŉ�^��D�a�c��?�9�)��.u[����mm��=n���=n�㶶q[۸�q�N���*nK��r[��e�[V�Ց�^�-��V-n��Ln{��rK!�r;w۫�Ց[�Ց[��u�[�8��g[m���q�r���E�[��Bܺ�m�qۅ�m9��n��n��`r[V�m&|��<<魎�R�m��sp&��������7x��Ot#+-��r+-��r[V�-+|�Y���|�x�A���ʭ�����R�-���n;��p�Vqk�VqK�m�[_�ń[9��_�V�ń�a�[L��L����f�m�n�ᶆpK��j��p[�U�[���	�*�׌b��;�+%1�y9�j�m��V�m��v���mi��Q%�}u � p;�v[�5�[ ���6��	ܚ��	ܚ��	܎��2����b��5�[��$���rok�Ձ[&����K9�mܖn �&p����o����o[
�m �j����j�m� n�߶�o�ڷm��ҾmE߶�������v n����}�־m߶�o�	����A�ȋ�@��%����o�/�v�m����C��]L�ńۦ�-��:����:���ۢ�m���m߶
o����x[ڷ�r�mǛ�9zp��D��w M��N�i�ݥ}�F�m}ݶ�n ��uy��Cj������m��#m�&p;�vk'b��mK�&b]����q]>�-���ĭB�*ĉ\��m�v �v��&N�R����*n���*n��l4?�3��ro���p�	�}ۊ�-9ܶ�m�V!n�V!n���E~ۊ�mE�D~"���O���"�m�߶�o�#�r���q���q���q[�-�ۺǭ{�"�-r܊ƭh���{��/N��}S�/n���*n��na�vl��n[���p���p��&p_��k�y�&p"W�}B��~ۊ�mE�D~� N�i{S��o"O��.ܚ�- �V�m�|o '򪺑e�[�����2��	�N��2�mE߶�o����- ��cy%|�W�m��D��7���&p[��5�[�5�[��~�¼- ��m� n��V�mk�� pێ��}[Ƿu|[ǷE{[��E{[���
��]���v�m����m��o"�j��V�m;��o[�7���
��Л�+�v�Co���ho+��K�������m��v���M����! ��- ���\�7�|�v��A&�e����mu�:p[���Vn��n}�p;Xy�'�}7�n��n��n���p�	��p+�rpk�&p����o���hok��n�w	ݖ�m�!O�/�8n�޶�m�޶M{yq�|"�� �K���m��V�m��V�mo�񶣉�m;�x�Ҷ.m[���0��e[^�mǛ�E�}[q�g����^�#B;"��8;���ߣ%��������ˎ��8���w�
|�
|�
|�kG�vtiGqvg��#/;��=��#/;��M���VG^v,�;����#/;���s�gǱ�G�vl�;"�#B;"��މ��`���A����Q�+��}|G�v�{DhGqv�{��;����Q���Q���D^B�W��l"?���G^v�eG^v�eG^v�eG^v,�;����Q��ٱ��X�wtiG�v��;v���D~��]�v4nG�v��;��#{;������w�uGw�q�־#�;6�qܱi�X�w�qGw�q��Gw�p��#�;�#�;�{�y�8�8}�8j�X�w�pG	w,ߛ���C7����V���^�؎w�qy,���#�;��<�[T�vtiG�vti�)�Ǯ��K;"�c1�	���q��D�ͧ^;R��H�#U��E��tiǑ�Ǯ��^;�c}�Q����tG�v�=$U������׎T��Uw�_{�_{�L{4nG�v�kG�v�jG�v�jG�v�jG�v�jG�vtiG�vtiG�vti�v�#U;���ڱ0�8��8M�؎wl�;���^;V�A�D.�;��wyx��׎�\��sy�>XmG�v��z�kG�v�jy���jG�v��;v���]u�A�G�v�jG�v�jg�Vk�ݱ��h܎��h܎��h܎��XrwmG�vtiG�vgyx��ұ���ˎ��8��X�w��_�D���Od�ٱ���{7�'��f{w�޻c�ݱ��(Ύ���ˎ�숽�]uG�u��;j�#�:ҫ#�::�c���Y+���H��S�먱���謎erǚ�#�:���<�0�ձ&�8V����u�	���W��r�~�c�ܱ_�迎��X9w�_G�u,�;����#Z��r�2��\���@Kv�c�~��%;��yّ�yّ�yٱr�(Ύ��X9w�e�����Bw��;�{=�c�ܑ�y�ђg�yّ�yٱr��ˎ���ˎ�s��Dhǡ�ǡ�Ǯ����M䱼�UwtiG�v�7�D^o0�{=�{=굣^�g�����-tG�vDh���K;���<Go�g���z�׎zm"?ѿڎz��&r��7���t�b���#{;��#U��u�׎�s�	���c��Q���Q�ڱ9��Ҏ.��ҎerGKv�cǡ�G%v��;��#	;��#	;6�I�{��erG�u�^G�u,�;����:ʮ��:���P�csܱ&�Xwd\�	�G�u�]�N���D_,�;�v� �H�nGvڍl�q��q�뱡���v�d���l�#/;�#/;���Q�[Վ�^��ؽv,Z;��֎jG�v,G;����qj��]ڱ�X�6��p��Ҏ`�`'��>�m�V�c�ڱU��ގ��تvlU��E�W��/"��(��*�&�=�ki���]����]��^��N亸�\U�D�C��8�*��m"O�[����'�^�Z�v�r{�r{Uu��������Dn��+���cqS�V�]�ݕ�]	ݕ�]��u���]�ݮ#m���ꮄ�J�&���WBw%t���WUwUu������]��q��ׇ�Л�+!ڻ6�]���]�^��^��y��r�~��@ޫ	�����5�	^���^��&�j�&�:����&�j�&�j��|'r��\��u���^M��^M������^M�D^{oi���2�+�j��p��p�k�� ^��^����:��:�w".��yׁ�W&xe�W&xe�W�w�~W�w�»j��㻖�]G�^�ߵ
�:}�Z�w��.��\�&�
 '���'��v��	���v�]��u��U^k��Lp"�@9x��צ�k��^1�U^{ﮘp"����^K�:���{w��Wx5�����	���k�ݵ��:��:��:���	����	'r���KF�Z���ka�U!^�V�ڡ7��r�۴w�W�8�� �h�M{W�x�{��{��{�W�x��N߽"�kE�uF�B^E�U4N�'�:�������0�
��z�Z��U�6�]���*^��|���|�:��:������:�����}���:�w"?ѻ�`�:�w"�OVy�	��^��_^��_^��o"�=g{�L^��^�D^	_D�7���d�"�Ǽ^g_��D.��.����+���^�UG^���#���{�)�D\�_��L^��D��嵵�Z�w�׊����ʉ���AVy-��k�ߵ��Z�w�W0y-ߛ�cy�ܢJ�k�޵C�ڡw|�»z�+����]K���*-���j(��vׁ�WVye���ג��8m���
&���������������{wu��޻�{���k�&^{��q�|�Z�w�r{��W�xe��b�kݵr�j'���4���!��&p".�L����i�Lp"֥������+�V�]g�^+�����ch� �
 � ��U7���泘����j��������Uw�ί�2��	��+���]�u�쵅����f���J���tW�w�9{�}W�wu|׮���:�k}ݵ��J����J���u�i�W x�W�w�~W�w-��6�]��d�]uW x�~W�w�~���4���k�U^��_�:`��	����	�&�j�5qך�k'ܵ�*�r�:s�j��pW&x5�Wx�~W�7���+�_ x�W x�W x{�����{7Q^��ut�r�	'��8�������	�r�Z97���+�}©�W9xe�W&x5�Wx�}����ʷm���]ߵ���BwE{�2�+ǻ�/�r�+ǻr�+ǻr��\�;�ʹ���_n�?�{B��K�]��RU���tj
�RU���t:�D.�͗ڻ�ޥ]u��K��R{7�׋���Ք�/�xi}]j�R{�L��ó�S{��ޥ�w��K�^:i5E{y�|�Ni_J�ҩ�)�K�^:|5�xy,����X'�����UM	]J�&b]��Х�n����nd�\��R��ܥ%w)hK�Z�U��BMG�N�9�:�R����T-��K�D���Ѯ���.Eh�tԉ<!�}�ʹԒ��l"/�;MK��˥p,�cis\
�R8�±��5q�%K��R^�򲔗M�U��p,�ǚ�cM+��ʹT����7Eh)BKZZ9�����-g�8K�Y��R^��cM��&��)���b�ԥ��\S�����\�w��D��G��vi�]��R��R���.�k�ؔ���v�T���t�k
��A�)hKA[:�5-�KA[Z�7�KЖ���¼�0/�p�K��Ot׊�R��_MZ*�Rq��ޥ�,g)/KyY
��F���p,m�KIXJ�R��ޥJ,%a)	K��R%�*�T��J,-�K��&r����R8�*�T��%w)K�X
�R86�w�D|��w�%K�X��Rٕ6ڥ�+e\�l�Tv��+5[)�J�V��Rz�Nm����*���䚖ܥ�+-�KWʸR��j��<�[t�E�[T��N�M�V:6m�KWZ����+-�K�W�&��؎7��l����]�¼tjkڡ�Z�Ԓ�S[Ӧ����p,�c)K�X���Z����^��T��J,Ub�l״i/Ubi�^Z��6�p,�c�״�/�c���Ԓ��l"��ĩ��%K��R^6���Fq����0Eh)B����!B����w Z�헎U���]��"��0m L]Z���R��0-�K[�R���T���{�KKZ�Ǘ��ԥ�}|i�^���>���/��V��.�p��K�[Z䗶���}i_�Ǘ��}|yB~�Pե}|�oV��/�x)�K9^:'6zi�_Z䗢��ho">Q��r���E~ik_*�Ҋ�ttl���9�)�K�^::6u|��K_��RǗ:���/��K�_��R�j�T������K�_���1���tmZ
�N�MM`jS���� 0�{�u�	LM`jS��t2m
 �n���&0��K`Z䗚���&p">Q&�2�t�m*S9��M1a�	SL�����/5��z�L��M�`Z����	�L0e��	LM`j�1�)LM`j�ɴ�d��� 0�LM`�&�j��0�) L�¦�]Ӻ�t�k:�55�) L`��R�j�����/�})���ˏB/z�ؔ�u��tN�D\	��RǗ6 f� �K9^:'6-�K��D��m����{�3gS�v���/�}iE_����ik_ZїΜMM`�ڗN�M�`Z�2��<��m+��>��|/m�K�`��J�W�ޕBo"�!�'��(9^�������z��+߼a�Tvm��J�W:���o"��̲0�t|��+_9Ҷi[:�R��kK�W
�R��j���ޕ�x%�+��J{WΜ-�ɖUxe^�{W�ޕh�D{%ڛ�O�Ѯ��+9^Y_Wr����vՕ�t�ڲ��t|e�\Y&W�-�^��J�W
��L�D{e�\�/WҾ����s%�+��J�W�˕�i�~�����q��+�_���2�r�l	 �ѱ��+k�J�W�-����we�[��J�W�{-U]��JUW��Е=n��+G����$t����r���ʩ�%�+q\��JW⸲ǭ�r��v���J/W�]k\��6�������w��+U]Y W��-�]	�&��ۋ������]�Wr��㕕se�\���~�R�B��xe]9��x%�+��N䱼�XLW�M��} �#mˮ� � �l�+M`iKX�����te�\�W�r�m��VҾ����~%��k�MA�W:�R�#mK�W
�� �,���Ex��:�+Gږ��t|��+�^��V:��8!;�J�Wv���+�J Xj��ڭt|���Ҿ����r[j�R��Ek��+��J X�r�mI�&��)8���[��rnY W��R��n��O(K9X���L�d�%,M`	 �!���+i_���j����D{%�+ߖh�D{�����p%�+�^�	Wvh�D{%�+��B�l{+��&���E{e�[��J�WV���n�,ܒ���v+�]i�������v+��B��w������~�Ȏ�-��J�W��-9^9���xeM\Y7��񕎯�w�����5q%�+��5qeM\i�J{Wڻ�ޕЮ,�+�]i�J{WB�r�mi�JUW��Е^��r���˕ere�\9�v"���Z�\��JW�����u����~�ҥ�.�l�+̖Tm"�Q�V6Ǖ�g�8+�er�K+]Z��J�V"�R���l"/�o�Z����c�ѱe�\�	Wv���d�%+�X9M��[*�r(lY&WZ���sb�ʹҒ����[�˕��[��R���q���c��ՒU�����$l"�����[v�p��RvM�	�Z%К�E�E�W%�*�JTUr-���myx���m%�*������*�Uٽ6�����<�Rc��,m+��D.·Z�����q+eW)�J�U���ث�c+����r�k��&�ǡ��S��G��m�+IX9��q+�X�������C���^K%V*�R���\'��!K�J�U���<!� �{-�XYW±R��J������!	+�WY�Vb�{��W�N�{������6��m���w�m��D����b�{M�{	[z5���?M�{	[��j��^M�i�aڢ�h�@�Z-�j瞶@�Zm�Z[��2��q����^kW[�6�v���Od?N���=m��-	k�چ���p���±���#���چ����mhk��!�-	kIX[�֎/m���kIXK����m�[�&r|Gnk�ښ��&�g�Ӷ&�Eh-BkZ+�Z^��v|i[&׊�V���-���O���˵�g�8k�Y+�Zqֶе�K[��"�V�M�O����-�k���b����m�k[������쭝h�J�����sm�\+�Z	��˵8��qyB�]��r����s�6d�\K��ʹv�i�/7������8��q��k�[�ډ��qk�Z/�'��kA[�	׎/m�Z����ms�D��o�8k�Y�	�"���M�'*�Z^���p�����V�M�'��!BkZ��Z�6���[�⬝��NGmZk�ZK�±�L��d�r������m��D~�{�ʹ����kZ�/זɵ�Eh-BkZ��ZK�±��5qmM�D~��֒��p-/kyY��Z^��ĵ���d�0�֒����Ow��Zq֎	��O�Qn�\��Z��"�V��@�ʹ֥M�	���ʹ�r���k-Y���1�-kg���r-kg�����d��vLh+�ڮ����EhmW]��ڮ�v
i����������j��щX���-���M����z������#hk��Z�ֶеz��j-Uk+��ʹ�_�m-hkǗ��t-h��E�g�[�Uײ������k��ڮ�VµsO[7�����v-�k	]K��x�:޿�vm�]�ZUת��˵^��k�\�&���Uu�����M�%�е����k���*��
��x-�kK�ڒ���n"�m��nr���X�y��<�ڵ�u-�k	]�Uת��е��%tm�\�/���е�X�b��<mo
r��޵���w������㺑-���޶L�u|��k�^�ע�v�k���~���s-��uy��n"��_Et|-�k;�Z�7�����:���5q-�ki_K�Z����p-�ki_;�u"'�OX �Ҿ�<��	k�Z��N�m` �2� � ���k�_���ѱ��k���2��9��&�2��	�Lp"?ї��Z����p�	lM`[ ך�v(l��N����qk�`+[9�V�M���`�[��6�W�?F�[_8�'�@Lض����m{k��Zr8���;�pm�D�����mab[��*������&ۖɵ
�-�k�ڶ��L�5��.�`�[&؎{m�`[9�b¶r����/l[�Z_��˵�c'���'����
�Vε�����T�Vε��0������ń-l���2��\��C�������m�k}a��~�n��*�v2m�B�XE��6�j�?D���]�4��/��\��M�E���0��v�����/j�ߗ�y��;��\��M�E.��Ma���ċ��ߗ�y�߯/����^���&������~x��r��w����;���п7����|�?�߻ɋ�q��:^�"~_�_�~o
/���(�{�
�"��F�=����{7�����<�
�"�����"Oۛ`r"o
�����w��+�{|����W������\��_���+��O�@;ދ\��^�~�>��uy7�/��cy��*����	�������y�`��\�wt�\�7D�8mD�8!D�8!��8G��D�s�7D㋸˻	��E�ޗ���D_��/�����a"���/�X�_^��u���"����E�K�݄��/�z���E.���/r��� &_�R}����E~��t�<G�t����{� L��K�������E|"Ct_�'R��"NV�"?������9�=i�"�	�~y��U��s�C�ߋ\�_X����E~�w&����O��ќ�o:L~���#�_䱼Q�"��[��/����|��˻	D�E^�9������ 9_�'z�a��\����X��E�6��E,��"V��h9��<���c��\�7�拼��� 9_�R}��v��E�}�6�yx�9p�y��M��/r~k�'p"�&���c�n� }���
}�'��
�E~�߇��/�'��'�yx��0(�E\�拸�~מ���T�拸�x̉�����+��qq��/���9�'�\�[C�"W�k��E.Ս��|��p#�9�"?�?l &_�'��q�/��nQ:_�	�Z���ȍL����D�� &_�i���T����)o
���0�"Αf�qx�D~�~��C�"Α����@Y�<����D�(>|���k-�y����E�S�'����y,� �ʉ�� �|�ڛ�|'����yx�+�#'�@ዼ8���;�{����4|Ǣ��E,�8�i��<��1}�O�4@�����B��c�����"��bX�\�Od`⋼�n+j_�R��"#m_��o�X��_����jM3��D7��E��m&��mEu��<�OQ�����G
_�" �/��`�q�宥��E�P��1�/��nQ���e��\�{��"�ѿ�_�'�`��E����̜�țŇ/��>k�k��Q�/r�ndZ_���G&��/r�nw0�<m��4��û�;_a}����'r?B�^�Um�(��E~��h��kB���<�ۊ��/���E���u��m7&�E��w_j_�"ܢ�&�"��i�׾�E��ۗf�	_�"���ȟ�_�i�"���������/��O@_��)4���7��~�ק����r�S~L̝�������r�j�E~"� ���j�E�#w�O&��?f��c��'�r�4��k_亸L�"�|�#�ȫ�v�(>|��go�}�����r�"�/�y�yHj��f�񉢽O��1��E,B��1��E~�F����>ߧ��$t�/r]<k?z_�i���v=��V�	�>��'���v=�/��������>�ݧ���w=�/r�<�>�ܧ���r�8��}�O	�1�v�?6ߑ?q�GO��������}�O�Q�7��"���N�擪}���<��&]�G�ދ\=o��T퓪}4���E��M�ܢ�O��Q��"?�?=}R�O��)�>Z�^�i��Eh��c��<���ӥ}��O����>y�'/��e`'�ɸ��CS�}4�ȥ��c�p죏�E.�7Q��^�"����"����±�9�yS�}��O�I�>�¾ȥ��%a�$�ct�\�/�b��������>��'���]yq|dʸ>��G�ދ\�Y��1��|2�O��	�>��^�"��Z����c��)ߛȽ-��4[���^}�v}���Yg�Q��"���Y}��OT�1��E^U�}�՛�-J�ދ��q?j�>��^�i��R�\�
�E~��ZJ�&r?2��E�N�EEUqB:�Og�Q��"/��h�{����Lދ8G��&r�2��E\h�֧����:��*�y,��2�O��1��E~��]��	�>��'���{���\���h�"���誛���Sc}j�Og�1��E����v?>���{�����6��F}r}��b�ڨO��I�>��Gs܋\�V��'q����".���S=M�?t?J�>��'q���{���~�F}Tν�����F}Lm}�?!��
�>��D~�;M��>��^�?���T�(m{�-^��Km/��o��O��&�}>R�6�;-�i�c}��w[Q��"Oۯ�����O��i�c}���]mԧz�TO���8}4�����0���E^/�i�P}�W��H�ڋ�9��S=}T�M�F�F}T���E�ݵQ��c��8|y�h�E��J�ڋ�i�>��&��*���Pyx�����3}t�M�#S��)�>Z�^����R�S*}������V��ї�"���X�K}i/��+q�$N���8}Lm}���{-�j/r]nw汾�O�1�k/��˥>��'�����"�E�D�4ӽ�"?����^ĕPc}j�Oz��&�}Sh��c{����Oۋ<���}�rʮ�j����;�@�h}̉}��;����F}ԱM�}B��I�����g����"B�m*�^����T����Q�TO�
��~?qi���iٗ�TOK�4��`#/��R=�l�%�ZB�%���+�v��u���j_�'rX��Ű��yyX�}��oΒ^-��bX��D�'��jɥ&�X��/Q�RP-�ɾ�O��a鬖ul�:�e۲{m	��d_�x�_L�}��ț�D~"w�e��xy��sTv-��N�CƵ0;�{[���P[V�-+ԖjKٵ�]KƵ� �"~h2�%�Z2�e���x�.��D.�]+�Z2�%�Z2�e��D�G����2���Z�%�Zj�eUٲ�l1��E����Zj���Zv�-��b��X��gKƵ,4[ʮe��Z>�=[�v}WB��K[*�e�ڲ/mY����"�}�V�����&�w [Ֆ�mY����"��=G��Dh�r�e���-�ز�l鿖%dK�5? ��W��*[*�%	[6�-��D��迖�kY/����O�^l1��E~�[�.��[*��[*�� ���qlY/��[b�eq��-��f���n+ƽ����z�%[��-��b�닼���`_�O�w �Ŗ�bK��
;��	]�ҥ-FǾȋ����cK��ti���4�y�~�^l�ҖmY��eK^���"N�q�/��X��;��aKq��[�-��R�-���mY��eK^���"/�߷g���\��]��tiK��ti���Ÿ����Z��R�-���\_��'z��mA�bj닼�nd汾�s���mY�mK�6�mޖ�%U[������.]�ҥ-F�N��.�%B��û�Eh�z�"�e���-��R�-[m���X_�"�OX�l	[LZ}���p��Җ-aK������û�m	[�eKز%l��l	[��%h[��-A��-+���m10�E����tԉ|�[��do��/�'t���8n1V�E�����miܖ�^�f�%{[���q[��q[�%U[vv-�ڲ�k10�E���6sO_�"|�3
�E~�{���<�_��{�"��~d��\���'�e_KU���"��[����[�=�ȧ��nI薄nI�V�k�[���ԉ|sW�-枾���(��-��&�� �[B�e	�b����n�to��$tKB��r���DӉ��v�-�Ė�ni�Vz�qlicKh�TuKB�l[6�-���-KȖ�n��	{ɖo���P_�'zSP�-{ɖho��&r�`t|ˎ�%�[Ҿ�\��!kϖ�gK�4��ڳň��.����/�ЖMhK_�,G[��� ����}�r��B\r}�����W[Ֆ0qY����K��Ą��/r~ɐ.}�	.����O�F&�4�K 8��+>Ѿ�%�[Ҿ%�[Ҿ%�[�-��b`�<��]���P[�[G���wKB��K[��-��D�me��R�-kϖ�g�Q�/�}S��lYU��*[��eU���-߲�l�������[j���[LZ}���C ���ڳ����/t|a�YXhj�P���/�}!��E�j�P���/�}!�i_H��r��-�� � 0�a�Z8�5d�!M` C v���X�y��	��B&�h��&�y���k�����0�! �_8i5lh`��6��L0�! i_H�&����S[�N��.�����x�;�©�a�[�	���։\�w��-���U�B92����nd�` C � �3T�Ҷ��-��BK�¹���� �my%x���mai[(���	�&04��	M`hC8�	�L0���� .�! `��B�:�P�er!���B����h/���ʹ��D� V΅�s!����Qn�\�/�˅&0��`X&9��B98���K�D~�7��7���er����!����,��(&��hî��/�|q"֥h����C��P�cX��ޅ�1�!_�bh'�Y)Ò�9��wa�]�{RȐB�2��a;^�#C�ȐB��WC6텵z��udH!C
RȐB�2��:�W�w&[�BC��L��1�����}!���?�ۣ�2�!��������K�R��U�ua�_(-ú�����1C�9[���}�A�����BVNZ�eh(��a��D��u��=f�1C|��_��r"Oȍ,���c�'e8C5d�!���B0��L�`2ԑ����:2��!�K�R���/ԑ����O<nQ'������KC|�ˉ\�_�l�e�/��pDk� z̉�D�͉�D_D$�!��C�V�j3T����e�/Þ��'0$�au�D��oB�plh;�{��s"���Jrϐ{��3�!�mgh;���pl�=�	���'���3����Y��]C�rω�DoC����`C':щ��JGC:
а1�G�C:���6���D^B_W,>'���^���P��Ň!0�i�I'r�:�a=bX�v!N�"ܢ�аq"�� �C���cF��$�a�aH4C���h�Ňa�a�6���Pm�j3�����c�3��!���ûz��Ň���f؅��3�����C�͐hN�%���`�z�Pm���!�!g8M6��a�bX��*�4�U�g9C��(��3�����fH4C�z�(o
��P�2� ���=����{Ec�����*F���!_�bX��Ő/�|1���� ����pNlؾΉ�c��zİ1�G�c�����=��c�zĐB���ab؅v!��2ԑ��udH!�Jð�00�Ȱ�0�a�a&C0�;@{��0,>�Ci��-�a�aH4C|��ho��_�chC�z��c�s"?���j3,Q!g9C�B�rN�|Ű�1T����fH4C�͐h�D3,d��͛�Vmn��s;�v�1��ۙ�[|�ŗ[|���[V�5�[C�5�yB�blY�D���-���O�>1���w�m!�_n��r�*��o���[i9�W�o'���[i���[i���[i������m!��cn=涐q;w"��}b�1�s�1���[��%��BƉX��r+-��[i��h�J���mm�v��VZnk������mG�D���-���6n=��cn�嶶q[ȸ����ŗ[|�ŗ[|�ŗ���<l�����Nߝ�c�����&ǭ��69n��Vmn���q�6�js�6�js�1�s�1���[i��Z܂�m=�Bn)�9nE㶆p�9�u�[�E��Q�[��ۉ�[���4���m��*n��v��&na�V!n��na��p�r�m9���-_�ZŭU�Z����m��&na�&na�V!n�V!n}�n1�q�	�&p;wk�&p � p ��o���Bo+���n�o�r�-�ۖn9�V�m;'����du�:p��^n+��mkܶ�m��&�X>�m۞�-h���KնTm[��L��j[���	ܖN��}{ԥM�?�UQ��Eh[q�m ��stÈ�&�z� ��o[�0��k[���j���^�굉\�/���mO�v�햽mA��mG�N�'�`U�m����mڶu�a�[�g[q��e[^��e[^�V�-ܖn]��m���m�n�ؖ�mI�D~������*���ح�N�ݒ�-	ے����ȥ���]ۙ��ѱ�־-�ڎ�ݖ�m��n���lm���@k�Ƿ5[[��5[ۊ���^ld�N��b�����ݚ�-���-������6�mk���j+��3g��j"���Fm!�Bm!�V=m��n�ӶCoۡ��Л��v�Y�����:���ڎ����m5�Vcm[���k'r�nd����}yxw�E~[����v�m���E~[8��c�.��V�Mĵw���o;Ww�˶u[^��e�.��g[q�g���-B�"��@��@ޭK�Vn�ږ�m��D~�����8ۊ��\��"�mu���mK��l+ζ��[q��	�"�-B�"�-�±-�Vn{�=��R���*�m��D,�"���ⱼ)�Ƿ��ۖ�m�ضVo[��-��±m��v�m���?!��V�mIؖ�mIض�n�Ķ$l+���k;w�U���2�mWݶ�n˸��k[_��][ٵe\y��ڬ��2���D{��k˸&���m��h��a(��v�m5�Vcm�ն�nK���d��j˥��u�T_�EU[T���ۢ��>��ǜ�j"/�[TT5����Q.��P����zڪ�mW�D��-�nQm�v��D��'�6��c?�&�=��K�ԑK{�%wǒ�#�:6���K��ꈪ���XLwTOG�tTOG�t�JG�tdIǡ�G�t�v;��u�Q'�u�QM�'�`=�=��c�۱��8�����訋��訋�`���H��p��cܱ ���v4HG�tG��j�,i"�Nst���8�������X w,�;��P�#%:N�=V���D~"�#%����ǽ)��ǽ��q���ϱ��(��"�(��"�(��"����jG�s��z�?Ǣ�c�ڱh�8i�H���U#��3m��{�z,m;��cC�q�건툗�x��#�O<G�t�Lǆ�7ċȍ�g:z�cCۑ8��?F�޽-�:B�#�zs^���>��q;r�#�:��G�Qձ��8:����\�X�v�R�Ҷci۫�%�i��q��/�ұ	툗�Mh�A��r�c9�Q=�ӑ8�ӱ���^vTOG�t�*;���z:�����W�b�9�ݭ*;ڨcUّK�Ŏ���8vDUGTu�ztVGgul;6���q�^�Ց^�ŎS[��c�z����f����hǎ�b��W��[�]b������8i��v�XG�u��zZ���q�Ŏ��ȸ�]bG�u�]G�� �����:�{=��#	;����:2���:ҫc�رq쨱����%���m�i�m;�#�z���Z�z�c���+�G�u,;2�#�:ҫ�-��u�N.�:j���:vv��h5ֱ��H��S�����u��:�#�:�cgױ��X�u,�:2�c�q��q�ֱT���@�X�uZG�5�Ku����uYGTu��zl�::���:�j���Y˫�sO�CN'r��u�֫��:��c��l����WG�ul�:NG=NG�ȥ���ꈽ���Xqu��z�_G�u,�:aM�9�-;*��\�ߑUbGv$aGv$aGv$aǞ�#�:���:j���:ҫ��:�P=VomԱz�H���P��[G�t�LG�4��w�:0�虎x�(��R�س5��wצ�����(�#^:�e벎��(��R�h����X^uGGptGy�>2�:�Y��Q*�ұ��X^u�KG�t�KǊ�#^:N!=V\��qr�/�ґ%�q���j".��WG�4/V���V��#K:��#K:6UM�'��,�:J�#K:�Kۥ�,�Ȓ�,�Ȓ�,�X8udI�.�DeIqx��&�X��#K:VIM�|�9U��u�K�*��g��O��;h󈗎URG�t��:z�c#ԑ8�vN�'��LG�t�:�F��,�Ȓ�,�X�t�J���c��D^�?:��8��虎��虎,���t�J���ͣg�⥫T�J��T�J�+K��8][����
����:Bs"?��~eI��֫g�θ�z��g��8]+������t�P�y�Wum^�B��z����z��,]�ӕ8M�9�E�J���کt�QWu�Y����z���k�ҵS�ږt�L���g�z�k�ҕ%]Yҵ@�Z�thy�T����,]Z^��U*]���x銗��HW�tUy�LW�t�K�j���'�+q���g�z��g��E��˫z�V#]��U=]�^^�^^���0��JWTuEUWAuT�T7�JWAu-P���v.�KM�"ܵ
����
�k�U]Q�U]Q�u8�u8�D�އ���ꬮ���u�y��r���Y]�e^�յ7ꪱ�URW�u�Wױ�Wgu��y�WWguuVWAuT�©��D�DUW.u�r�+��vP]յpꊪ����Au�vP]5�Uc]Gh^����0�TW�u{y{y���2��<��!eוq]��hM�i{�q]��h]�K^���l]5֕^]�Օ^]���Y]GB^GB^5�Uc]5֕^]�?^�?^5�UcM�����+��ҫ+��ҫ���
��<�[�"����:��ǫ���W~[�&b]h�ҫ�\�� a]�ֵ�:��:�q"��w ��{]��u��T늪��ꊪ���:��ڳ5�W½-����+���j]������zu�W���?e]+�&�}
���UqBڨ���ڨ����^]!Ե���Tum��r�+��U���zܵ�^]��u��Uc���׺���D_�e\W�u5[W�u�ƺ��P�+��ҫ+��a]յ��*���������&����5�յ��:��J��EXWzu-ºj�k7�Uc]���EX�"�� īٺvc]5�Uc]����k"��Fh]5�Uc]5��Y]벮uYW�u�XyB�Z5ֵz�^���g�m\yx_�-�2�+�2��ٺ���ٺ���ٺ6{]�ֵ��ʸ���ʸ�f�
��m\�q���k���l]����[W�u�ޚ���]q��]�i�W�u�ٺ�e]벮J�ĮJ�Z�u-պ6h]�صA�jɮ��Z�u-º�+/�±k��Ւ]I�D�C�l���^]-�Ւ]����l"������K����K��l]��u��T�Z�um����ޮ������^���u%tW/w�qW	w�pW�v-�J��q��kAו�]�ە�]�۵����u����Hȫ������}]˾���ꮃ#���ꮪ�:Kr"Oۛ��`�J�����������[ކ�9�?o0v�]��u$�D��/"Ҿ+�6�]Ǯ �����J����J����:%��%vu|�z�+�Ҿ��N��Ҿ�<�7���  ������]i�u$���]��u��u��U�]��U�]�ʮUeW�7o�^o
ҾkU�U�]�ˮ��ZUv��x�~W�w�}W�w�}�Ɏ�Ɏ�1�W x��a��ڳ�d�kU��^M�u�� ^��R ��T���/����,mK`
 S �j�T�M�	�#���� N��O�&0�=K�`��Ɏ�ǉ<�=�=�ȋ�kA:g1-G�����!5�i9Z:g1-GK��R9����r0��i�Y
 S �� �Mh�	L��&�4�q��i{Y�^�2��	�&0m/K�_���	�yB�G�t��D~���s�)ӡ�)&L��RL�����,������0ń�L�`�ӡ������NG/��0?���05��	LM`jӢ���&0-ZK[�r�>��V��X�ss�u>ńiC[*S&�2���&05��	LM`*�R������h)�K9^:�1z)�K��R�7���;�}ii_ZJ�Rڗ:���/�KK��R�7�W�[��/�~i�Z
 �
� �C(S ��teJ�RǗ���h/E{)�K�D�B/�c��cy�㥭ji_�D�G�B/z)�K[�R�����o"��[T{�ڻt$dڄ�
�T�B/z�Л�m|+O�^��R{�6��'S��6�M���r�ڻ��,�8K�R��n"�=KK�]�q�r����+'�n����}i�.�θL`:�r"�MA�� � 0�) L��R�j���-�vK���j���-��}a�S_8���ED��*Ĵ�--mK}a�SL���tgZږN�L1a�	�Ҷt�f����t^f������#9L��R_��X��0ń�p��r0�) ��cqq���K�_����t8f��&��a�~iC[:/3-mK�`�ӆ���-�^KGh��k�����0ń)&L1a:{s"O�ͧ/L}a�S_�V���1S�j��X� 0��_�_ڽ�� N�O�Ҷ�	�&05��.��2��	���	LM`jS�� N�R��N�L�`��2��	��/u|)�K9^:h3�x)�Kgo�j��K�^:/s"?�-*�K_^�I�Жj�����/�}i�[J���i�[:B3�) L`:B3���� � 0�) L�_Z&��ɥ&05��͔	�L0e��	LM�D~�w&Gh��ryx�L��M�"���S_���T�&0�) ���{JoCj�����/u|��K�]j����M���)��+�&��7�^*�R��
�T�o"?��.Ǜ�r��U�ڻ�ޥ�.�v)�KU�D~�{[h�N��s��B�>�Л��U9^
�&�⸑�w��K��Rh���L��D�ro��Z��0/�r��ΔХC;�¼�<Go
ڻ��e{S�ޥ�.�w�hω�D������nw��Rh� M�]Z���M;�R��r�tLh��RU� M���.�vi;^J�RB��Mg���.�v�д�/��K�]:4�w��K�]j�R{�ڻ�ޥ�{��K����DS����}|)Ǜ��sS(�^9_�D{%�+�^��ʊ��~�%�+��J�Wr���M�{�J{7�L~"�e�D^	n
��+�]Y�Wr����zek_Y�W�/-�D~"���t|e�_I�J�W�����t|%�+��J�W���h�D{e�_9�t"O�[G	 K X������t|e`9��,,���&��	,{˹�%&,1�|�y�({K&X���\=o�,�`�&X/"�,'��cUK_8���=���R!N���B,bYVX�É�D^j&����JÉ��ކ�%_,�b}��
�T�e�a	K�XV����U,�b�	˂����%&,1a�	KLX6�̈́ea�K_Xb²'��	,G��Ձ��ֲ:��,ab	K�X�Ĳ:�$��/,}a�	�R� � ��}%�+i_��Wj�������{Z����t|��+��ʊ���M��P�ܦ��X��z%ڛ�c�~o�^9C��~��+�����	���%��E�Em�+M`i'�J�������p��	'���G`	 K X��}|�t� ��Q�>� � ���Z����&�4�eE_iKX�FvjY�W����گ�}��P���}ek_��J�W������+i_����|�z��+�]��ʁ�����ޕЮTu�X�r�ji�J{Wڻ��l ,��J�W�U-�^� 8����R����y���`�~e�`m�'4��	,M`�&X2��N�'����i�ٮ�lײ����Z���X����Z��R�r�l&,1aY0X�r�d�� ײ:�Ą�,ǽ�Ձeu`IKr8���c��D^	�&�Ē�sbK_X�²���%&,1aYVX��:nw�a�LX�-�
'�X~1P�5�e�`�9Xb�rl9��Z�v-�뺷U��B��E�� L,ab�K�X*�R!�
�,+,�a9'�T���ز�p"?�Ec)K�XVN������R4�|��%_,����R4���ea����R4����[��rl9�D�%L��MA�Xv�0�T��B,�ɖ0��,b�K�X��$��K_X������,i�D~��Q�W����e)`I��i�eu`YX�-i_I�������~e`	 K X��U�� � �t|e_ٴWj�rXm	 �a�e_��7��Ѝ�,�`Y�W���8�r�*K&X2���	Y�WV�� ��}%�+k�&r]>��_[��i�4��	,��&��nwߖM{e�^Y�WҾ������Л�O�o�:�R�Bo"W﮵�l�+i_Y�WҾ���h�|[v蕎�t|e�^I�J�7����oN��u�m9��z��+�]i�JhWV����+{�J�W
��ޕ%we�]��J{Wڻ�ޕ���ve�]9嶬�+��J�W
�r��D޽-�+ߖSnK{Wڻ�ޕ��l�+��J�W�h���[v蕎�E{��k9�D��t+�Z���՝����6�o��kߖ� ����k���Z��V�u|m�^��Z�ע�����w��k��D�8���?�9m�^k�Z{��굣v�Z���M�"xso�^��Z�ע��B�z���ݤz��k�^����ͽ�r�����n�^[��N�mU]�ZU]��Z/�J��i��p-{k�[��Z�ֲ��i��p-{k�[k�Z��R����<��Q�-Bk;�Z����w[���V��z���R����T�-�k��¼�X�ƭ�۲���8굶
o"��V��R�����jq	ui�ۖ��Tm�?���cWێ׺�vXmK��޻���T�����m��D��V�[k�Z����Ѯ5n�w��u-�k%\+�Z��ίm%\+�Z��vյ�0�굉��_�z�Ķ.�ui�Kk�ɶ.�uimW]��&��rݺ�v�l;M��k-U��c�|���%wm�][r�vյ]umW]K�ڮ���n"W��ӥ�.�ui�4�v�lK��F�V��m"�+��v�^k�D,B�ֶе-tm�\�Z��"���f�2��L�-�k��Z�֖ɵ5q�^kk�Z��R�������^mC[�Z��b��ǭ�^��jeW˸�ѱ��j�V[�֚��ڭe\m�[os2��l�f��kW;s�e\-㚈u)�Z�՚��lM��}j�Z��V��k"���j��Y���EU-�j�����ǭ��:�ǿ���ZA�v���km��D^h��q[��ZTբ����uVmC[�&�}�Y��ҫ�^�=n-�j�UK�Zz�:���D�j�W-�j;�Z��j�vtl����Vc���O����>!�j5V��ZT��ĵ5q��j;��9�-�jU;|�m{k��ڶ�B���P�zjK��Ҷ������B�����QmC[k�Z�ڨ�F���P-�j��Z�ڨ�F��m����F�6j"?�]�>��KkQU��ھ��Y����Kk��ZTբ�N��d_Zۗ֎Um��Z�ڨ�	����r��K��Q[A�NGmG��j��j'��ĩ-Gk�Sۄ�z��	�mBk�S��Z������UOm9Zۄ�6���mBk��&��⩍j��Z�B�V=��D�ڳV=��gm�Y�&��E�RmZ˥Z.�v��6j"O�ǯ��-GkG��Mh-�jQU���r��	��R-�j��ZA�r��	�T�>~�Pm�Yk�Z�N!m���SH�&���8<W�&��Ь�/��Fv�hK�&�X�mHgՎm�UK�Zg�6��Mh��Vc���K��E���l�f�Zm9Z�Z���h�@�Zm_Z[�֖��f�5[�`Ҷ/�5[��j5V�Zg�:��	m���~Q�gF��]��7�-����\�������ׂy%~�#��O��O����}xQ����E��0��������E^��;��\��M�E�����"��{x���}yx�������"/���Ë\���ċ\��}�E�����"�����"���ׂ������\���E^��{΋\��=�E���u�E����q%�P����E���E��
��zoV_}�'����E.����E.��Jl�ߗ�y�~_j^�/ g/r]��+/��Yф�"?���W_��_D^���:^���`�^�'z�@����孃ڳ���K�"����ց8{����A�ڝ�>��".�k/�	��"�z�E~�7�^�"����6�w\ڋ��_��`�jyS�����o�E.��ً<���'^�p�#�&r�#�^�'�Z�%�Ƚ�%{��woc�^�"������?Y��u���c{��(3T_�?�OCۋX=��E.���ۋ<�[��"~�c{�W§;ul/r� m�턩�/���|���>� �^���vB�ۋ<G��p/r�<���"�B�"����E^	oC��yx�d��^�'zϡ n"o0@�y��MPu�Ca_�Ue�8G8ދ�DoCL�}���C'܋�Do0t½����E.�[��E^/�'�v/�W��y,o�U}���nB�ۋ�^~� ��O�>��țh�E������� �{�'�k�j/���T�l�6Ek/�A{/��r}�_�� |��r�S��"��q�S��"���Lp"�;=n/�X�mL�D�<P��"?�o`��s�@ۋ������L�"��� �"?�7�&�B|���M��"/�7�ľ�O�>�B|�W�7
�^�/��!��<m�9X�q,���9_���*�d��T���	_�R�O�_�	y7����n&|����9�"��; ul/��x�h�E�>Ek/r��m��D�6f_�'�g�<����}������������E�6��E�� |����r��M�����".N��y�/��|���_����(m{���!�|����Hۋ�^~����E�k!�/rnd��D�Z����E��F!������B|��w�S��"�ч4=n/����G4��K�h|'�h�ȇ4|�E~�/�����O�r|���ց{|?!z�^���e�:��z_���"W����"?ѽ�B|��w#_��!�U|��-
9|���-Z>~!�/r��DF����c�	_�R��:���"��V�{�E�+rp"��9}��Ї!&�E\{ ��\�o�h��� ��st�10u"7 �E~����"/���ػy,��R��"�哏
��r?җ�"���S��^�"xi�(G{��'~��O�7��">Z�^�"x�~����EpS��P{����	�E�;�' ��j/���.�W��/�OL��)|2�O&��?��D~"_�?i�D����G�ڋ<<�џ���}r�O����>��G9ڋ<Gn���S�}�OB���>�����`����7�Oh7��woK�>*�^�	�g�O/���>拾ȋ��>	ݧ���rcB_����T���ûk�r�^���}L�|���y~�^	���S�}J�O	�1��E.�W�V��w�}t���E��eo���O����"�%���p�I_�i+�&�I������|����"��|��^�'z��m"�|���������������Tu���[����K_���鮪�$tul/�X�m拾�c���r�^�[�!��{�E\/��G�ڋ<��ZA�'h��kSH_�i3�t"�@�1��E���}��M�e��<!�����}�}�?4���������FV�}t½�u�ݕp�p/���v��}9}�Ǜ���Ӹ}4ǽ�O�M��y��'m�z�S�}굏��yq|��>����O�}�O��Q�"�f{P�}�����/�X����>:�^ąf|�D��w ]���щ�ی}��w#��>*�^�"�#�GM�D>��ey,���9�E.��ۊ��i�/���e&�D~�}�O��Q&�"~���.�ӥ}��Oq�)�>Z�^�	��&r]�<P_7�o
�O��Qr�"?��{�ۧq�h�{�����c��\�wf���+��¼������0�E�W~A�Gaދ<�� ��O��I�>��G��D>ݥj�.m"��D��Q�7���٧8��Uz��}���/b��M�}�)�/���{7�{�F��z��p죅�E��;M%�QL�"~���"��棫�E^	��tս�O��K��	�"O�-ʴ���v�ҡ7�/�O��]_�ui�y/���er�D>�)�{�K�/n�_���{�"�J��D�Z�^�Rui�v���k�z퓪}R�O����>]ڧK���{���M�޻y,��K�>J�^����t]�'B�g���S�}��M���}"�O��)�&r��S�7�۝��/r]>��k�z�S�}4�����N���O��Q�7�߷gqqDh��Vo"�v���e���C�E����{���՚¼yx���6M{/�}`��\�OwA�'h��r���>]�'B�(�{��w#�{�"��mE�݋<���޻y	��i���ɡ��}�O���{7���*�q�m_��U�}R�����|����E\{拾�M�Dn+-�G�܋<G������|�2&�E��_bui-t/r���B�"��G&cB'r?R&�"W��S��'U����"��-k▖liɖpl1{�E��X±�[��-���r���ڥ%��c���l"O���b��<���%[V�-y��Ƿ�%[±e'ܲ�mI�kYǶ�c[��J��^K쵔]KƵd\�
���D���/��&�Tb��ɷ��"�[*�e�ڲ{mY�6��w#[Ƕ$a˾�%�Z��-m�ȋ�~�xd.�j�ȥ�%aK���K[��e��R�-I�D.����x�.�q��s�{�hmiɖ�jKK��d�q�/�y�.���-��R�-�і$lIMhK���_K���^ˎ���8b�e��Rv-;ΖgK���^�9�/�X��9��]�5���Y+�Zʮ�\�۝����e\˾���8�K��KƵ��"���Vٵ�K[b�ń��.7��jK�$a�ڳe{�{M�"ܢ��%	[��|��	m"?�ǯ$l�q���"?�-��Z��p�ɸ��e���e{�{-גq-�ʖ�ki��fki���j�K��XK���X�^���Zj�e��U-�Ė]b����G�%�Z6�-ǖk����bK�5���x��-�Z�e	��l-���l-��h-�Ŗ�b�ў/�n�;@_�R��6�-F{N�@�d\�Ʊ��Zʮ��Z2�e��Rv-�D�h}"��-a�J��<�Od��h-˾�e_K���WKz��WKz�tV��%�Zҫeq�D,B�5��8li���`�J�%�Z����Z��\jY��TKA�TK����"?��hK�b�苼�nQ�Բ8l)���a�.7��j"���J���Zr�%�Zڨe%زl���DU˲�e��U-˾��ji���^�f��\�۝��/��L!}'t�X��,�Z����h-��h-��b��<��m�ֲ%l"O���k1��E.�o�w��;�$l"�=G%�Tb��9±�[��e	ٲ�l����j���L�"����V�M��o�L!}����ܖ��\�Ow5֒^M��J��-a���/��E�WKz��WKz�l	�����Zj���Z�M�'��Wc-5�Rc-��&�}�3��E�N(��K'r�����k�%�d\�+�_Ƶd\�.�����o
2�%�Z����Zj���Zj��ƚ���� �uX/��]Kٵ��D�tg��D�ZK��ZK���[V�-��h-枾�Gy�`�D>���"ᭃ�/r�Md\K���g��cK��4[K��4[������P~鷪l鿖�k�K�$aK����"��}��/���^���:�{[%�Tb���/�}yP�-k�&�ziɖ�liɖ�hK^���"Α��y�Bm"OȻI{7�UmIՖTm��	��-�ז.m��v�-�і�hKж�j�&��8[����yB�mƗ��ûkgKq�gKq�,G[���8[�e�b���5ao�MÉ�a�Y(�&���{�BqZ�pViXU����,�d�`�p0i��BK6���5=�e�%-Yh�BKZ�pV���(Wv\׶m^a�E�"�_�+�g'f�߁���Yv��}�]����F�;rh/�e!���B�h�f!�v#'�Bg!�m!q�e��,$�B�,T��Z��Z�%�d!�Bh!������KV{�xٍ����U���F^	6ð�3T��՞��,l�Q��K���K��PUg!q��n��]��e7rx����/K;Æ��KJ�B�,$�B�,����/�P�e7b���B�,��B�,t���#�#/W��Y���xY���xٍ�U+^��B�,��xٍ��W�,t��Z(:C-t����!�g!K�da�fؽ�e�%,��+4C�,d�¾�/Y�1{�PBJ�B�,$�BUY�*���K���Kz�B.-���^�y�n�ri!�z�BT-����ZH���Z��ⰐK+4C.-�����ri!�*�¾̰/�F��[�z�{]b!�bo!���n����{�6��+��.�J�B�-��V�1��Z���z�B;.C�,ԋ�z�/]b!^�ew9��>4���ȱܑm��P��ː8�/���ŧ8,��B.�FN�MZ�X���y�e�B�X��E��K���ڍ<!7|k/C%XH������Bh!�Bh��+��B�,t���P�Bh!�Bh!qgaUe��Z���,YȒ��X�8�d!8J�B$�F��%*8��B�֍�Ю4�����d�T+D�B�V(�
����
����
����
a�г�]!�2[!�Z!�Z!��8�4V�Y��UHP�ȱ�˗Xm\�z+�BW��
�[�z+���[a%d��
=[!J�B�+�B�+To���г"a�z+��BJ,��BAWh�
)����	�$CgW���(Kj�B�W���f���2�����K��P�g!K�d!"a!�_!��]aqd�q��?t!�q�-�!�v6�n���
�X�+��B+��B+��B+��B+tc�n�1�͎aAcHc�4VHc�4VX�4�4VHc�����
�X�+�B�*�B�*$�B�V�+M֍�^n��?���!�rV7�1�'䪵�1�j�PUU�PUU�UHP���a�c�F�lTH=��S��
A��z��(�P!�P7b��Q!�f(��L!�z�Bx)��B�V�3�<S�%��#�:4h���zu#����Q�>���1Ē�ǐT�q��1�B�(4U�(Qh�J���JK�RŴT1�R�Uڠ��حR�(�W�tэ�^��g�2Hi]⍜���.J�Ui7b� ��k�+e�%����*%�ҺĴ.1-B��CIj�J��KJ颔.JQ���F~B��Ԡ��D�T+���"�9{(S]V��JI�ԍ��K)���K)���K)���J�.+�e��R�%�XR�%�����e��#��"N)�V/�6��ƕڸR6*e��6ƔzJ��TЕ
�RAW
B� T*�JA��JkS6*e�n似��J٨TЕ
�RAWJP�lԍ�^��lTj�Jm\)A�
�R�*ťn�$���F���zJ���A1��R�Vj�J��\.wA�qڲQ)�V/�Ջ�\ۋ��z1Uo��TZ���R��+%�R6*��n�i��K=��Rj�JuY�.+E��ŴA1��n�]i6(��)��P7�\i�R�)��R�֍���L)����R7VJ*�XR�%��yD�U�`d�n�X�bI�4SR)�KL�^��Ǖ&����R�(�%L�8J���.J�S7V��n��J!�J�X)7���Rn(�^�DP��JW)7t#f���E)]���R�(uc�n�K���r�k�J�SVJ*��R�z��R�)�n�	yH� J�R6*mPL���TJZ�������Q
�(QZK��E)7�rC)7�����%J��JW��*U\��)p�Z�R)�^�XR�%���i�`J*��y��� �R� ��Q
�֫�AJ��AJ��AJ�W7�?� �R�����XR�JI�Tq��K)���J��*%�RR)�^��R�%�>��gu#?G���rqJ�qJ�X�+uc�lT
B��SZK�Z���Oh���Gt���J�W7�*�RO)��
�R�T
B� Tj�J٨�.��P�p*mL�qJ��]0��R�)�����J;S*uc�lT��JEX�+ťR\*ťR\�F�'wq��JZ)��PiSa�F� T
B�<S�3��R
/��R
/��Rj�JZ)ϔJ�R]V�8��S�g��� �}u^��Y�����0�%LA���0�R�)��R�U�J}V��*5U�����J	�9��V�*%�R�*ťn�|,�T��Ri�`�K��1U���J����0ťR6*UI� �}���~UI�*��JA��J�R)��RO���F�UK�j�R6*uP��T8��Q��*uP�UJP�v���J٨���F��Y\*ť���p�R)g�BU)T�ڥR�*�n���P�$*�D݈k?n���U�Jq��p0e�ReS�F�ȱ�Ƿ���qՊ^����p0-Lѫ�]0��R#Tj�J9�9U�4�MiI`*cJq���ÿS��R[\j�KmK�Ֆ���R[�Ӎ<"�[�j+vڢW[�jUm����ikq��R[\j�Fm٨-�U6mA���i�Fm٨��i�gڂP[�Vƴ�ܲQ[�ҍ����m�J[��F΋�����-��-	܂P[�i�3my�-ϴ�1m�-�E�n�9~�V[?��ϴm�RO[�iK*��ٳ�mI���iK*m{���V�噶<�^��K[RiK*m��-]t#���7�⸐冶�~[Hh	m�J[nh�m!�-$�u*m���Si	m!�q%(mQ�-������^��m��-볕m�G[�э�^�>[�gۼ���j�-س�_ruF�j�-ųmEE��-سmY�-�{�:�m5�^�H�e}�ң-�s#'�6'�e}�5{[5�Vz��muF[�g�3�A["hk%����A[w����û[Im����-$�%��D���-�%��Dж�oK���]�A[+���?[�gkښ���z[���BB[�Ж���mY���g��lY�m���ٲ>[�g�l)�q�x�ϖ��";[d�F�����w7��R<[g��t�I�l�D[+��J��m}C[�Ж��R<7��~��7}YL׶��Vg���t!� ��?�����GY��6h�p�%��D��n�Aۆ�-�%��`ϖ⹑û?���8[!Ж���9[gK�l;�L�������s#>Z��|ΖϹ���Ldgkڶ�m��-��5	m��-��5	ma��hK��ȩ�:Dc�h̖��r0[GЖ�����z�����H��i��6�m�@[f+��/۶B�9	ף ͍��;� ͖��
����--��e��̖���2[4f��lA�9	L�\(���M����ųu�l�9�+M�d˛ly��xg+�يw���Tيw��ʖ]�R)[�ΖJ�R)7�Z�-�r#���OPe�l�<7�Gq���gK���I���`n�$\���.-��e����$��m�yDN�e��>a�ۍ<�w����h��l1�-f��l�h�����mK�n���I�f���hn��257�z	�l���h��Um1�9�7EE[QѶ6n���x���p�Ev�0�}t,�9�������*���o[�fK�lɛ��h�la�-y�%on�	�L.y�%o���VT�ۅ�>��3��S�_XDvv�B,y�%o��h�.ں��0��ْ7[�f��l���j�q��mۖ��ꌶ���p��x��l[dg��l��yB�ㆯ-iK�lJ[�g[�-q�R<[��V���x�j��i�ضU#m�i�{���-�S�=%�S�=%�SR<7��e*)��Ϲ������MIޔ:�RgT�9���$oJ���A+k�J��djn��ޗ�MIޔ�MY�V�7���,8+D%�S��tJ�P��K^25%SS4�6����L�ƔLi�)ј�)јRTz}J�O�ƔhL����KI���J	����yD���])�:�?�$\J΍��\Cr0%S�wJ�N�ƔJ�����^�ְ�p)58%�r#����)9��[�F�K4�F\	�n�$djn����Z���.�����s�R���)����)�<���t�.���))���)���ͬDvJcO��)]<e�Y	��ƞ�ͬ���9{׶DPI�DP�fV
�JH�$�J�O		��P)*!��TBB%TA�#��O{�FN�{�(Q��(Q)*�B�\��Jਤ�ʲ��,�,K+�D%�TG���T��h%�TZ�J,�d�ʲ��]TG%pTG%pT�D����#�Ln�Z� �RY�V���k��,^+y��g*+�Jĩd�J���6�RT���D�mI���l3+ᥲͬ��JQQ	/=���<ӓ�q�RO����J���SI=��k%�T����S�3*�D����J���V���*�D%�TROϨA�K*��A*uF�Ψ,K+uFe�Y	/�V����y%�Xm3+��RATG%pT��J�P)*��K*��JR��=B���]CRO���ѽF�����S)*�Be��挜�/�֠���C\�<G��%��@��Az��H�f(�����ȱ|��T:�JG�������Q6�d�J6�d�JGPY�V:�J\�d�J6�d�JGP�K�-k�I轖9	�G}C%�U�X%�U�X%�U��J����J+�{.0rx�L�JQQIc�4VIc�i���MD�ޥ0r>G� *}C%�Uv��ȱ|��$T��r��*a�R.T�_%�u#��;�V����d�Jp�F�K�Q��V�e%KV�d7bǧ�/+���pT�JJ��b+)����n"^V�e%^V�e7r^ޙ$�J�d�J���+;�Jp��J$�T#�W��e�ʎ��*ѫ�*ѫ�*k�J�Qi8*����*�J�Q�q�ң�#����V	h�ң��*���I��n��h�\iK*1��*��*��*�Je�\	h�N���*ѫ��D�J��D������*	�����o��J���JR�$�JGP�*��JmPI*��j%�T��n�i�8��SY�V��n��}&��*��n�T]0��J��>�8�;߸��F����~B�|T%AUT%AUJ�����z�\�F?�r��$����J�QIP�t%.U�Q7��|��ʾ�y��t*��I�8��R�t����ԍ~�W'q� �����>l{D6���F��F:2[Gf�F�_7��I�FN��xt*1�#�ud���֍�+�q1�c�ܑ�:��a��f��[��r7�X�G��Q�t(JG$�{k㎶���{�HGҍ�����pt4G�^�#�u�u;�^7r.Q��c��іt�%Y�#Kv�%��y�pz(�n�G�r��Q�H��K�c�=mGz�H�Q�#�vD���MA.�l�����yS�q;���q;���۱\�F^�ܱI�(�:RuG��H���#Uw#��3�����.u�厼ܑ�;�rG�XTw$�$ܑ�;boG��H��c��Q8u�׎©#�v,�;:��@ۍ�><,�����ڑ^;����ڱ����#�v�W��#�v�Ў�#qv#�w�J������F�W�cGJ�F��H��.u俎d�Q8ul�;�_G��������{�p�W8ul�;�]G��Hv�QG��{a�#�ul�;�^�V���pY�l��cQݑ�:���ȫ�z����AuDEuG����tY�^ѫcGܑ�:BUG��(v:Z�n�ݚ��%n�ƶ#ud��lԑ�:�QG6�B���]0���������YURGo��u��N��4B���#����:��URGf��7w���r�r����蠺���fh+�Q^u�WMUGJ�H�MU�:�#Kv#&!^vT\���$�gG�����cQݑ%;�dGp�H�uYGJ�h�:�cǢ�#Kvǎ��#%vtcWG��;*���ؑ;V�+莊�9���
�#qv���tG��F?��z�j�ˎx�/;�dGp��:Rb7b��_G��{a�q������:2[Gf��l��c��Ѡu4hѫ�����ۯ��#guT\�ߎձ��HPK܎Ց�:���%nG]֑�:TG��H=y�#�t䙎��^�_Lᥣ��%WG�ՑT:����iGyՑT:BB7��_y�>��&TG��Q%u$��D�Q%uTI���7��:�EG�Աx�X�v�T;2HGo��u��tэ~���貒:꟎(�%:�����#Jt$���ϑ�9���`�ٹ_)��S�F��7CJ7��ۉN�#�st*Y�c���9֠JG�ѱ�������r)hK:����б���}�S�t#����ѱ���fvl3;�JG5�8:�DG��H��#�s�����9ڒ�DБ:";Ǟ�cOّ�9�9�R�#�s,%;z���Q�t{��#�sd}��ϑ�9�>G[ҍ�e���F�e5>�	���#�s�%���@�؟vd}Z�Q�fւ=-�s���hY�������E�e}�γ9	�c���ʦ�����?����Z֧�8��O۲�Am�Z	��#��[�S۲ֶ���Q�(Q�c�m���i�V�����P	�'2��}h��yq�k[����Z����Z�T��m-��:�Z�T� �ҍ8!T-��bI7��k�j�T�����Zx���Zx��Y�<S�3��RK�]l-JԢD-J�rC-�s#/!;r�����iY�9�k[�FN��涱�49U׶�nm�[���N�0N���I��U\��N��j����i����i�U�\�R<-��
�����.��9-�Ӫ�Z>�UI�*���i��ƹ�Gtc�u#O��(yӒ7�$��l�ڸ���4�ũmk1�V�Ԛ�Z��gk9�����%�����imI--�ֳ��L[��4-@�4--�6��������G��Զ׭�u�p�H޴�m-f�b6-f�25m�[�Yjɛ֩�:�Z�RK޴�͍<!t�ln���2�kɛ��i�K-y�:�n��X��ij�Z�R�Yjk�Z��(�`O�Tj��֖�µ�p��%�n��}Ɣj���j���j���j���j���B��j���iJm�[���";-����Ӗ��9�.+ɛ��iɛ��i������c��hZ��hZ��hZ��`Z�R��֢1�y��^Z�(݈+�@�EcZ��`n��.+ј�iј9	�D5/�楶���lڢ���i+��
��i��i�V��25--�ʘZZ��3�Mr-S�25-S�Z�Z̦hZ?Ӎ^�Rk^j5Km+]�Yj[�Z���G�K7r�Z��,�|NK޴�MK�t�Ь-��%�t�-��%��N�촶��ή(��#���U#��΍��K�|���r�ZT�J�Zd�5����pԂ=7���p�Z�Z��-�k�����U��Okj���$�J|Z>��k���iU?���F��&��";-S��ｘM����+�c��MK޴�M[��
�Z!P�����i�?���FN&�ӂ=-��6����1�`O[�֪~n�X�iֳ�������?m[��i���j���j[�Z"��xZ���qZ=O[��";m�Y��i���i��칑û�T��O��i����EvZd�Evn�}Y�iMBmZK�ڠVԲ>-�s#�ruH�O[�ւ=-��֠��g�ק�<k�>���%�Z"�{Z��EvZ̦���ȩ���L����e�x�Ev�R��i]<-��R<-���yZ��EvZ=ύ��5�؇F�X�v��'4֠�DЈ��������������yڬ�칑G�l���`���Y��)�����n��aՎ����|���|�h�����3�F�g{F����6�>#�3�>7r�Mn�$������7�>7�Bs7�I�F�O�#�3R<�oh�������}s#�3�?#�3�=c�HތMr�6�FN��Ց�ɛ�1���3�ˍz�����Fc�h���F�g{F�g�xFc�h��;�RgDvF>g�sF>g�sF>gT�J���)��[�F��0���ȱܷ����q��e%�3�7c��h�a�ьs#g�՟3�8#y3�q�����m����џ3�>#�3Zvn�T]��?#�3�wF��F��ۯ�Ш�����m���^�џs߶<!��z�1U-;c=��]l#J4BB�eg�Fnh�F�g{F�glF)�����F���)�ь3";#�3";c3�H�����lDvFYΈ�����|΍ޕ�4����:#�3�>7r^�G���xF�g,K��������F�gd}����Y�I~���G��WHh��FHh���j#74V��(э����t�H�t�H�(�X�v#'�mHi�F�� �r�yD߷��Uo#�4�Lc!�(�B7rx���74ʅF�it�<��3����46ɍ<��3݈#�8���h��?c��B��ӈ8�Mr�h��Ӎ��l�loRO��g��F�iD�F�id�����A����K��Su�Z.7:�F�il��9��
�F�iD�n��>)B� ԍ���t����gAc��H=���h��q�q�QA4RO#�4Z�Fj��l��FM�g��h�q�QAt#Oۇq�����zEE7����F+�h%{�n�'�@w��.�n�7�7
q��A��K�F�illuF#5�P��h���.��z[��J�Qg4�F�шK������h��ң��m,^ѫ�ѫQ�4��F�j�O��S�w ѫ9{�9�9/W�4�Hc��ٻ�ml1���Q�4���4ֈ^�N�у4rVc��HP�j��?mڕ�i�n�iK=��Ӵ_r��F��h8uF7r,��퓨 ��Sv#��O��&.u#'�Rh���HPM�%׃t#'�7ڲ������z�QT4V�� ԌO��n�-^٨��=H�i$�F�j� ����F�l�(=k�n�9�\(u#��G%k�f��H�j(�P�hK�H7rx׶��ƚq!�Ai����ûD�%:nM�X3�RJc����Y��Qz4J�������E��2
�4�FǨ����f�"O�諾��%�"'�w�ȱ�>*�����_�T�>=�����"?����F�Ջ<��e�"���z�_��O�/r���w/�z�]C/r^�Ћ�8w�9տos/r���9����"O����������ߍ��2��U��"�<Ӌ�=ҋ~�W�#
�q�X�n�w�}�S�����#��Q�~F����y^�pmCP��#���<{�'�w�}������yB�:`�^��O@=�ȋ�w�}��^���B�"�ꭃ�y뀠z������E����"��>A�؋�=�Ӌ�CD/�;��>��Ku#a/�����"g��@.�">4�B/r�n�`I/r���/�1���AT��X=ǿ�Լ�y�}=}�W�y�Җˊְy��yя#z%�ݡ�^�i�Di {�Su�BP��[?7|��9��6Ջ�=2�9��W�1/��9��/Ս�����:�{�ӫ�]� N/r^.QZ�^�T]���^�R�]�"��	�"�y�.>ب9	W�Ӌ<G7C��^�9����������Q/��/=e/r,��e/b��J�zz5�N�g_@�9	�_<H7�R�E�ޅ���E��},�EN§Z�yD�L�y�\��?/r,��t�O��6$�"�w����ȱ\i�?/bx�1��(`ϋ�����E\/��q��?/r�4��9��_t_�p=��"'����q�Q#��r�Fg�"�w�8z��w�ݮZ��y�]۠D7r�cKz���	��yD�;j�yB.w<H/rx��z�ϋ�A/��+�ϋ<�?*����]�ы����ENµ��"�хL�؋<G�6ң9�_��E��p����˧m��n�&��"��%
��"O�Ň��E~�Ei {����
�s�!*zя��كټ�#�ټ��]C�5��"�|΋�8�8/r^�!țy��y�E��w\C�9/r.+����0�9/��~B>����r��ټȋ��y�Su)�{&���C��$�">4�A/b��27r)��{�B/r����}.�7�">4J�^�\C��^�܇�^�\Vt���J<H/r����{��"�ѥ y�"'�>DOً<�?�`8z�G���ы��|T�y��p��k�J�����K�Ћ��q�A7�s|���^���'(�ȱ�(��s�>1�'��^似O@�ȩ��B�ȩz� 8z�G�I���y��2�-n�E�˻	tы�>ՎO� G/r^ކ(q{�W��D����΄�E?��i{��"��n�I*}2H���'p�	}��^�w�����8b�yD�&��҇��E�[�G�ۋ<!n
���'��8}T���Ǽ�<b|�P�p/r�<u|إn�oVިy�܆>�Q/��}�^�y��p=��+�}⓳���>q��Ӌ���Q��"�����ĥ>q�O\꓍�d�>A��z�q��8���XN���O��q�D�>��� ��I=}RO7�C��)�F}�n�r�z���>��oԋ<!^2>��^�	���n�$x���F��#��ť>�Q7r!K=}x�^�$��?�P7⇳O�飱�E~�.��Oۋ�^�Q�����Z�!�������'.u#���F�"�w��Y}rV��Շ7�EN���oԋ<"/���Շ��F�4q�9U�����T�d�>�O�F^	7�傑.��z{eӋ�=~�9�����1/���Ӎ\0�	L�:�8��#�%�x�E^/��b{я#�e�g��>y�?Ӌ�>v�3����t$�>��O,�x�E���eӍ���3��#��	/}(�^�$\��L�n/��T�$�>�N/b�X�n�c��҇��E�6'��!cz�Gt!�%}��^��r�C��"O�Oy�O��^���>��ҋ���	��/�O���T���#zS����cyS��(�{���.*.�!P�?c}4ɽ�Ix�������~�9UoȘ^���Q6��#"cz��gzG��ĸ>��O@�C�t#�D�>ѫO��C���G�zy���D�>��^����^}X�^�����>i�O���;��/���gr\O/r�s$�>ɮO����$�>$Q/r^ެ�F�����������E^ho0�޽��}A�t>J�^���_���'���}x�n��DJ�	�;�����>��OJ����{�G��#��������Fp�C�"��ې,�'K�I�}Rb7�ކd�n��爗}�����>!�O�C8�"�&�� ���O0�j5{7�y���@�@�|x�^���U+��I�}��^�X.Q��O����"���'�����"�w�
�}Bh���� ��!�z���X�7�E����j��'q�a�z�Su�a�z�Su���t#��@ۇ�E~�����Iԋ��nҔ���"���D�>I�O���{�-��I���ٻ�ڝOz�^�D�>Q��^��Y��5���E?����V���E�އfLU/�.>��^�]��q�$�'	�!�z�ûD��>y�O8���څ,�	�}�q��-����z_rJo�wȫ^�i��}BhZ�9�[�\�'^�I�}����(%v#������EN���F�9	��\�'��ɥ}ri�\�'��	�}Bh֫y%�ȥ}ri�\�GSዜ�7Q�O.�C��"�� ��ɥ}x�^�$~����>���gk��Z2nK�m	�-�_�����ES፸�,Q�%��DՖ\�B[gK�lI�-)�%v��U�ֱ�q�X�dKAג%[�dKg�/[:��ή��kɒ-5^K���ٵ�|�Sem/��%q�$Ζ��Rе$Ζ��Rе$Ζxْ%[J���/�∗-�%^�t-m\K��B[����9<�Km	�-!�%��$Ζ�ْ8[gK�B����n�� �To-��%��$��/�B{�8[�eK��F^/n�%�>!��4{-�^7�����y���[�pKn)�ZT��y���n�T��ȸ-�_������$܍���%/w#��iyg��[RuK8n	�-�o��6�9U�:D�=�7�>��l��-�_�9� "U��-�f���yD~�X�wK�n�*����=GU٢z�F�MT�-�bKo��-q�%��d�n�cxf/��T�-��1	9�%�w#�^l�[r|K�o)[�}K�o��-Ѿ���Fх��l�.�d+��a�*���J��[zɖh��8��^|�c�`���8��[�Ŗz��^lI�-	�%��t�--a��q�4(��I��"���	�--aK�nI�-�_K�nQ^x#���pK�m)�Z2nK�mɸ-�%���Җ\ڢ��E~��9�;�f�9U���ڒ^[�kKTm��-Q��l	�-�%^�dɖ����k��-Y��l��-����kɒ݈�k��O>����0�_K�k���"�r�i㺑c�\(������ע��E^B�ĸ�׍�}HkIc-ѫ�gk�ٺ���%��ki�Z���ȱ\|Z�ʾ9Uף�֒�Z2[Kfk	h-�Eeߍ\|4�ȱ\��XKk	U-�[K�jIP-��^�$|Գ�$��Ւ�Z���st�U-��%Au#��.*A�$������u#/�w 	�%A�ĥ�����k	U-�_���IxP	v#���EZ7r^�e��"��>!ٵd�]/bxɮ%ٵ��{׋��9�w %dK�k�l-�a7�B���"g��ql�q-�bK�ؒ�Z�Ŗ���Z�^K��F�3�d�R/�$����R/��컑�Q�F����U�-UeKfk�l-���w�e%zu#>4i��>�*4[t��ȱ\C�˖��EI��<m���ZZKkIc-i�%��t�-�y��X5�-��E���<G�E����/�1������%��h|����W�k�q-j	o���Z�]K�ٍ�����%�u#��Jb\���1	:_�$4�-ɮq%$��^�%���-�_�wBJlI�-��%��-���%l���ȩ�eJv-ɮ%��D�����Z�WK�j�F-٨%u#��+m\iʾ�P��Zʾ��Ւ�ZrVK���ZBUaSa�F���!j�B�)4{�f��������
٨��0�x��ԍ�~ڡ�+$�B�Vhк���Jq����i�K�lTH=��R��
y��g��Sec��гz���
m\��+�3�C\*ĥ�/�!�Q��+,A��
�Z7�C�
q��
q�9	W�lT�F���:�n�U��
�^!TʾB�*��B�*��B�*ĥBWh�
m\!�z�B�)� �����P��+d�BWB� TB� TB� TB� TB���!!����,d�n�y �`7���+$�B�*$�b�� TBU!TBU!AT!AT!ATagc,�9�{��PB�R!.�R!.J�B\*t��lT�F�lT�F�z���
�c!�P!��B�)��B��Fѻ�Ջ��,��� T؍v#��T�K�u�!A
�n��� �Q!�P!�P�	-4��&�������C�*µ-TBU!AT!.�R!��BZhB�e�����kﲲz�F�Rh
�B�YHP�lT�F���wd�g!TBU!T
�"\�:�B�Y��:�B+��B�Yh�&�q�b\�-$�����
j�B-��B�+T���W�K�o�cx�ѭ\�ڍ<�w j!j�BJ,t�E�o���&�/����#qga�dH��ȱ�������B�%C-$�B_Z���Y������qg��,��B�,d�B	Y�%�e!^�ea�dh/���K2$�BUYl����\Zh��	��9U~sUe��,T��@[����!�m��,����[h/'C�-��B�-T���[h��9U׶�P/�k!�vI�z��^2d����h��h�c!�m�^�Fћ��ۍ��w��9]b�K,�ޢ\�2n�%,��B�-��B�-d�Bz-,��O�~�n��k��+��\Z���ٍ<�{�ZH���Y�kH�+t�]�!��_��+�x�HX���HX�ݗ&��	Y�+�5^!��^7rxwQ����"a!"a!��BJ,�B�+����	�^7�}h	��P�u#�r3�`�,��n�]�g7r.d]b!�Bh!^v����\������݈O[-��B-lռ�û���B.-��\Zȥ�\ZX���B%XȒ�,Y���X�^y#�ѕ&K�d7r>�j	-a!^�e!K��B�,l���	e_!ʾB�W����	��qqD��B�P���B�W�^�d!8VU�,YȒ����������2�K(�ʐ%'c`NC�,ԋ�z��%��B�,�����B��û�E�BT-D�B�׍�C�\Z��ZH����!�Bh!K?�1�[�z+���z�TЕڸR�Fg�:�RT-t��Z����I�I��yD�{
�����L��j��+m�L+!�J����k)��:�R.-��L5^��+�����ٕ�?�@[���ȱxhN��T��e)^v��w�w�8K��TЕ
�RAW�옲d7�]|��R�V���dWZ���X��*�RyUj���Gtu{�dWڠ��])ٕ2[)��Z��*�R�*��n�x�K�Q).��%��T�K�����sQ*�Jq���JA�qJy��gJy�T�6(�����t#�wkZnMRO�7�F�}�RŔgJy��T1-UL���zJ���TJ5K)p�G�S)�R�RZ�x#O�e��)��ʞ�9�ۉXR
�(Q�g�ëlJ�M)��bI)��bI)]��E)]���n�X�����Y���r�����~7ImIi�ajK����/�DP����OjKJmI)���>7rx����Rd'�%�ȱ�ދ��M�٤�MjKJmI)f�b6)fs#��\�&(e��%��1)�V	��Լ�4)-��2)��,)Β�)�.i#`�TJ9�zI�K)Β:�R�%%\R[RZ�w/��J_E�%�v�y/�YR5RJ���Jʮ��ʍ8��ҩ��,ie_�YJ[��2�zI	�Լ�.)Β��Rv%UR*%�RR�R
���J
���J
��TJJ��z)����R*%5/�Tʽ�8��rV�TJJ��N�TI���JI��Լ��*)��"()��"(�-)%IR5RZT��&7r��2����۽���'�r#�w˔JI�Լ�R))����R�R�Y���r��]��+)�r#�wm�gJ�L)��j���I�K7��(cJј�I�K�y�F^U]Q��j�n��֡�)u*��P��F\/�J)S�����#��3��z7�Ҽ��9)�s#�DOa��Iɛ�I1���I��n��Ф M�TJ�R�&�lR�&�lR��F^	��hR�&h�N��Iј�I-N��)Ec���I�K)s#�h5^�Ƥ�K*cJ�����e5^�����gI{�R�R
���Լ���RZ�FN�e%@��2)-�ʘRZ&�`R�F��F�R
���KjKJ9�Ԗ�ڒR4&�%��L���L*PJJ)-�:�Ҷ���I5K7b^4)-�r07���eRZ&�eRZ&�eRS�FJ�R[R�[�z)�
�R&�^R�R�����y�\�r07�]�r0i5^J������.�^R��F���]�%%\R�%%\R�%�,������I[�R4&Ec�̖��ʘ�h����,7r<�n��-o�� m=H[e��lmI[*e�7�u*��I��n��N��Si�lA�m�܍<"+mk^ڂ*[�ּ�5/mq��fiˮlٕ�Si�7�%\��r7r�l�[��T��c��>^<��-�u*m�J[fK�܈m��V��(mJ[[�֖�� m=H۾�-f�ej��6w#O�mn��lј-��^n�w�)*ڢ1[4f+*ڢ1[��V��`��z�����z�B/[��z����z�B/[=ϖ��WBfK�l	���g+��6�m	���g�l;�n�cx/�;��ˍ<�+Mf��٪~�g[�f����m�>7r,W�����z}�����b6{�D�l�L͖��J|�L͖��25[�fK�li�q�h��g[cύ����xg��l��yB�i�y�z�-f�-8����T��g����$��?n�@[!�����v��%��-kۖ�-7�mYۢD[�VA����l[�FN�'d�E�^�-���my���h�8m�-ⴕm����hBm�G[�і�ڲQ[�����ǻ�PՖ���n��m����h�Kmq��oh�Km���VT���n�$�ˉ^m�E;}w��nk%�BU�:��]���*��r�mw�V.����4֖���X[k�p�E��
�-z��mK�4�V�E�n�w��+hm}C�һ-Ƶ-��b\[Q��J�%��=x7−][�kKvmɮ-���m��-�u#�r��lm��-�u#/��+b\[�k+*ڒ][+���Z7��^���n�𾨫�я#�q��-��2[[@k[z�e���֖��Z[�Ж��2[7r�ZMB[�Жٺ�^fk[��5	ݯ�Gtm+�ʅ�5{[p�F�ޛ�,ٖ�Rb[+і�Z��H�	�Z��H�	��^[�k�qm�D[�k��b\[�k�l�ȩ��Ÿ�4֖�ڢW[���9�z���rV[��ޅ�U��h�Y��ƪ�h+*�rV[�jKPm}C[�iK=m�-�t#�ѯ���V������K�bI7������GXᥭ#h���L[�iK*���}�<~��{k㶵q7r^.y�m��V���n��~��Ӷ�nK=m����gK=���}����m��
����V�ť��c�5IPm	�-�e��l��$�m�ۚ���Ӷ�n��:��t7r^>�
Bm�@[6j�Fm��l�������V����<Ӗg��K[xi���L7�"N7b,��m����RO[�iK=m��-��������#h�ڲQ[6j�Fm٨�6h�F���ݑe����V����B�=>v�J�ťn����P����W��U9�9������rV[�j[��嬶r�-g�嬶�ն��QzDo
rV7�{qJ\�ĥJ\�ĥn�c�����'�һ��SBU��쮻�߫Z�X���F�B.��*�@%�U�W��D�J��D�J�Oi�)ѫ��z,A%zU�W%gUrV%gu#�������*�����$T��J���JGPIP�Eue+]�K��T�*[�J�P�*9��������+���*�D%gUrV%Tu#g��]t��{U�!�4�W�q����\��JwQ�q��V�l�ȋ��Z6ɕ����*;�J�Ѝ<!�K@�F��9%zU�W7�Jh%*��*ѫ�7T��J����J��7T��n��e��ⵒ�*��RTT2[������9����Ս���2-^+�҃T2[%�U��J���J@�T#��֍��7�1	��{���*��Jث���z��*a��*1��*��J��ĸ�J���*����*mI7�R�T
�J���'gUrV7r>�
U�PU�F��l%.UROe=[i^*ᥒT*I�K*���.*颲R���J�8*[�J�d�J�d�J�F��OI��T��ة,K+�N%�t#>!��K*��.*������t=���8��Gt��U�JR�$�JR�4B�ei�$��JR�ĒJ�4B�F�K*�9�[���R�t#O۵-�T2HeZYpVG�7�d���R%UG%pTڥJ�T�%�ei%�Tz��f�K*�Pe3Z	�tQ��g%JT����Ѝ�5$7T���n�*�M%�SZ�JeӍ�8>=�VA%TA7�n�A%TA%�S����T�>����J���J���xJ����Gt)�l*�L%fs#��L�$oJS)c*��ҼT���"��)��n��[�`OI�2�*�Q�T�=e)Y�@V֍����⹑��z,_{J��T#�mf%�S����O���mfe�Yi^*���*!�R�TʘJ��F����.�y��Ͼʘn�i���3��RY�V�L���,K+�����8��h���FN�_t-K+q������s���K��T�Kݥ�	�`Z�F�����t#�L>Z[�V����U	U�����*	�:>)U��#z��*+�J����J���T+�Q%.Uz�ną�*��J6��K݈-.u#�wmk������ AUT%.U
�J���K�v�����K��U�Y�©�x�tP��Ս��k[��tP��U�*T�p��b+ѫ�.UڥJ��F��B���G���D��z�q�Zec[	h��Vi�*i���*i���*T7������U�*9����tP�]l%zU:�JU	h��֍�^>�l��V�l��U�^��U��*��J@�������*��R�Ub\�.�l+�R�UZ%�U*�J@�*x%|,�*EX��h�:b\G@�X�vd���nG@���:�����yR8b\G��F?����<q����׍�7�����m\Gב�:v���cm�	;"a�ڸ�z�Hv�ߎ�#�u�l;���}v��Z7rxn
GJ숄�����H�������7w#O�6�tG���:j���ّ8;:��ڑ%��K����:�������!�#�v�Ў����|�M>�&ri�N�#�v�ҎmyG��Ȓ-a��>!^v����#qv�!��%�H�-aG�F���9</G�؍�8�d��u�鵣^���cG�ؑq��X�+܈�˸���X��e|G��;�Ŏ@�U;ri��#�vԋ�#�vDՎ��QvD�n�	�OGq�U;�jGT�ȥ�aGq�B;BhG��H���9	�r!�#qvd�n�\|�Ŏ�ٱ����w�ٻ��z��u���n�		��bG�ؑK��P�ؑ^;�kG�ر��(;��N�?��!�y�����Q�uDՎ������]GAבq;z��@�h;z�����g��o��n��kG.�ȥ;�\�Q�u�e�bp"W��Q�ul<�jG�֑^;�kG��h;mG]�h;겎}�G����#�vl*<겎�B{�mF^	׶�W�e�T]�ri���ȩ���ˎ򪣩�Ȓ=i��Su�%;ʫ�,ّ%;�cGp�)��\|vY�c��Q^udɎ,��yB.+�UGy�B;BhG�(�:Bh��f���֦£��	��<���Z�#���HFNU���Tx�ޞe��#����:겎��;"tG���I�#	w$�}�G����^^���y�#/wT\}V�>�c�ᑗ;�����#/w��}�G���gu�Tݑ�;*�����;�vG���F~h�Md�$�QquT\=���y�^�����y�#/w�厼ܑ�;�q�v�c���w�����G�����c��Q�ud܎��h;�����v�c��h;�kG�֑K{��F^�jeɎ�#8vǎ��Q�u��;�cG��;�c�^k�U��ǎH�Q�u�Ď%�Gp�Xxǎ��yD��ή#Kvd�n�9��ʒY���눗�
�����u#�*v�jZGJ�H��Z7�x��:J����;6Y�#%v� <v������p!k�:�cG�֑�:v=[7r.>a��T����#�uTo��#v�%<Rb�*����h�:�cGp�������ȒY�#KvdɎ,�Q�u��n�ܤ�}�#%v�x�]Gp��:�c7r�>m����#�uĸ�ב�:J���ձ]�U	�#Au$��"�c����]T֍�ЮZѫc����:�Ww/�;�VqղQ-��RO-�t��G[%�Z��v���j	���j���TjMUmI`K*��RK*�U����Z��U\��S�8�"��]��^� TK=��S��bI����Z�E�n�T٭Z��E�Z��E�Z�U[�w#NH���Zn��ZH���k���j���j��Z��e}Z-U����V8u#g��\�Amo`	��st��(э<m���Pk�j��VK�j�Z-Ս�Gؖ���m�E�n����?����}c�?�Ϫml��i}V-�ӂ=7r^��Z��A�V	��O����O��jY�yq\|Am�`K�`O��`ύ���Z��i��iY�V8u#���J�T���ȩ��V	�r)�j�R-�A�p������p�5U�Z��j������w!��j��iTmo`�������i�7��Y�>�������*��z�Gm�`� �n�8j�Xmo`��bI-��2H�T���F�ֳ�z�Z�e�Zਕj�R+�j��Z,�e�Z]V� ��э��n��Aj��%���]�z�Uo����>)h�jA��j�^j�^j�^j�V���L-���L���E�ZAWK=��Ix�R�ղQ-�Ԫ����V�����<S�7�[-��ROm#`��䪷Z�V[�ת�Z�֍�м)h�jm\-g�
�ZW�K���j��Z�V��j���jm\���-	l9�qUE�ZΪ�x���7rx�ήyD� Toף���j٨�jA��zj�^m�_[�ײQ-����ZR�%�ZR��}��m�_+�j��gjy�y�,Q�rA��jA��jA��jA��֖�%�-A�Tm�_U�U��ײQ-ՂP-�RO-��RO-��ROm�_/��].w�`-���,��"N������\��&-u#�r�B��7rx� �R-պ�Z�X�غ�Z%XU�U�K� TK=��Ӎ�7|A������Z\���U��j�_-g�*�Z��FN�[����Z�W�l��+�3��-�Ւ]���F�����V�l��V[��*�Z����dW۠ؒ]-����Z��ŸZ��Ÿڞ��֒]-��b\7bxi���j�_7bx�`7b�*�ڞŶg����	kK[qX����},�v#g�@���Zث��=��%�E�Z����m�-�*�n����'%�4��XK��J��k���j�����2[-��Z-���X-�բW-gu#�(g�rV-Tժ�Z�V��jq�9/�_	������r�Ԡ�T�A���Z����Z���W��9/����Z��-��9����U\�򪖠j�[�U�j[��� li��z5��FSՍ�Nul�U#�u���1�����i���p��F��h����b�1�����i���i�yD�k�±�p��ƒ�y�YV#�5��F��X882[�JjĸF�klUR�Jj$�n�,>����(�5�]�Jj�F�]��e�{���{�d׈q����]p�?�����4�_��ila��]p����������-N#�5Z#�5Z��iT6����l��֍��5j��n������z�G�Ӎ�!]Oc��������pD�ƊÑ�O��i��FJll=����p4B��#K6�d#86�c�$j�Fp�F�'�UR#86!�v��.5ڥƺıqD�FTmD�F.m��n��c]�X�8�k#�6��F�Xqx#�����H�����T5ri��j�R��ڈ��\�ȥ�>����X�'��FS�ȥ����T5�j��j��F-�����#�6ʫF�md�F�md�����ŔqGzmD�F�(�Q�U!�B�X7rx� ��FTmD�F.m�e�֫��q,{�W#q6Z�F�l�^�,�Ȓ���������H؈��H؈��H؍�hU\��؍�;�����͎7� 86�_#�5黻�����Su!��n���qa��#��e�F]ֈ����/Z#qv#��o��˵-q6g���F��w !��8����5��F�l�q�,�Ȓ�,�h��9/�g#K6�c#8v#����(�я#z��Q����k$�n��>��k��F�lt��(պ����}����F�l�l���H��R�Q�5g#q6�F�ld�FJl��F�k�F�k�F�k��F�k,�a�9	���'wK(GJ�FN½V��Ȓ�,�(�Y��%Y�)�э5�c�ktc�,�XBy#'�B�8��ѳ5�P��/�%�����j�����	���8r,��#G�ktc�d�X�8�]��j��F�kĸF�kĸF�ja�"���i���G@k�F@k��Fk��Ƃ�Q�5�F��F��g�㖩A�FN�_�4h����Y�P�ؠ8BU#T5BU�klP�W��j��F�Ս��ťF�HP��HP�ՈK��ԈK���kĥF\jĥną֠5�R#�4��Fxi�Y�>��q���"ı�pl=�yD70��g5�����QK5"N#�4�K�7j$�F#Ԉ%����]�F\h�P�j4B�<�(��Go�B� ��A8�Q7r��G	������±�p�F�j���9���pD�n�w!�A8v���l���#�5�F]�Hv�d׍�WJuY�k�F���l���Hc�4�@c=5�?��(�����O�����/r��w�9����"���ϋ<�߅�"����_��n�/j���E�w�}�����_4D���z��߽�E�������#��~_�	�]�O������"'�wm��I�ݷ_���_�����G���>��I��)�������?��1<H؋8G��yĿO
/r��o�/r��7��%�"�ѻ��݄��g��^�������Ix�A/�"���G�y��8{�'���E��߷�yBކ����f��"'���^�E��}�I!���P%�ԑ^{� ��K؋<���G?3%G�8{'�q�E\U ����==������"�=�������<զW8�"Oە�u#��֋<��c�:��������"��L�ߋ��߇��4ugz��p�D	v#��Ջ��kΪ��Y��k��E|�W/�J@c���"{�X'���z�G��:#�_����A=��/r^>�b�z�c�Ұq�ȋ��"��Kg׋���g׋��K��E��g�y	��Po�ȩ��Qo������"�r!CP�?�q�@U/b@U/b^�����I��A�"��2Ջ�Cta�^��>�"�z���� A�"���W�9	_��^�$���Y��#z뀳z�G��T��� ��E��7�yDww����ց��E��o���^�X���^���R/�T/�qD� ԋ<�˝>����zW��E^ߑ��^��>ZCP�ȩz���F>) U��K��F��4����T�"/�k�׳�{B>��Y��� ��E��w �_�	�|��E��7d_����X���Y����1�� �u#2�Ջ���^�U��z������Tu#_u�q��I��"�z�c�8�ԋ�^n�ظ^�9�j��X>��K��'wp�yD�1{���v+/�;�9���׍\�8�^��n�`\/r���^�X>ߣ��!��#R��"&q��)B|��E��[�׋�; �׋<!�r4^/�qD/�>,ً���
�e/r��s��(�yU�����_��>��z�Wջ	6��o����y��bPb/�qD?m��q���z�WL�a���zã�z�c��^��>����I����n��%�">mJ_�i�D)U|���8�/���g <[/�� �^�w�aк��6�9/����^��cz����׋��[9=�/r�t��"O�UKyዘ=\ڋ.�E�T�E�U���E?&�9�jA�^�$ܑA�^�$\۴��#����^��- z�F��; @ۋ��|?n�@h/��Xa�^��ZX��rM��<�����9����yD�6��9���@h/�|roí�^�D�>�_�w�@ۇ��F�`>�c/��M>Z"o�}�q�d�n���?Z"_c��s���>��Uً��x���>�%_��)|��^�$��?�_�$X�Ʊ9/V���U���}"a��/�D?��q؋����؇^�>2�D�>��Op���Gt�~<|�e��/�JH�}�e�,�'Kv�cyBlҟH�'��Iv}G���]i�+�.�����<��^��'�u?���������#���q}H�^��.��w�.�yBl�^�yD�x�^�٤?Y�{ً~L��/�d�>��Op����>)�qڂcB�q��MZ��/���{S@h��i���'��>�e7���K�"�r��^����ږK�����I�r�ɥ}(�^��<�(�^�]�X�^���(~w ���VT��EN�%*��	�}g���'^��{�Gt=J�}g��ٍ���4��9���kw��}���">G,a/�s��J�=G7|�`/�>`	{���//�	�}�p��9�7�_/r����!�z�Su×q�d�>�^7rm�}m7r^?ֶۯ@�'���8�"���E?�+f�>Z��x#��\�'q����"�r�O�8���>:_��!��O��ó�"��B��"���H�}1h��I��+��	{}��^��n�"a=�/bxɮO��F�%��a�z���$�>1���qqĸ>1��R�9/=�7r�Iv���]i�_���'����z���^+��	{��K誕���q��ȍ˝O�����>��O��C��"���]��C��"��r����>a�׋<�w ��O��.�EL�֋��b\_�DŸ>tY/�R��+��a�z�Gt-2m�7�V������>a��\��_��yD�Z��O����ĸ>1�O��F�Kl��˧��%V����EN��a��O$�	��x��_���>)�O����pv��I_ue�>����q%ĸ>i�O����$�>�[/r,�%�>	�9UW�P�'T��F}�P�/r^�4�o��EBU�P�'.�Q^�"?ZW�qY	U}x�^��.�
_��)���g�"fOy�8"���8"�K@�����>i�O�����>i��>����9�׋<���׋<G �Of���d�>����yh�q���#���^�E��7ѫO�ꓳ���p�m�t#����v�.�E�@f�F^h�����I�h-��*{�@U�">!a�O��A�E�˵�q�EN�p��Of���p����C@�F��k{\��X.�9�Y����"�壵��'��!�z�G��Z@���E��]�ꓳ��l|��r��^}T��'A��}����K�ג�Z4ވ߿�lԒ����Z�PK�i)�Z�PK�FΞŷĥ�J��l�F-�_�o�K\j�K-q�%����K�ע��E���ZrVK�������f�E%�<"���Z2[�J��I/�`K%ؒ�Zʾ��7⦰���dג�ZZK@k	h-�_�	�l-i���k	h-�%�����֒�Z�?��;��%���l-j_��]�rV7�;��kIc-]K@k)�ZZK�֢��E?��ٳ�.=[K�F�UK�㋼<4/9��zk	U-�_�ח}{IP-q�E��^\j�K-�o��zZ�8ވ�����Z�P���yD�#͎/rx^���U+u#�wmS�x#ףf�%A��}-e_K�j)�ZBUK�j	U��#����n�	���;�r!/�_9��%li	[Z�ՍK���ZBU7�uv-������n�T���yD׶բz�E����9��lԒ�Z�Ö ԍ�U+��䙖��%��-e_K��qZ�LKgגgZ�KK��R��To-y�%��$���ҒAZ�U�/���"�%��(|�Su)�;���Ҡ�����Ң]�EgZ�KK]֢��E�5$�t#���ROK]�R���� ��Z�P7�]|�RK��ҳ��l-�
o�.*��t-i���k	h-�%���3|���Cfk	h-]Kfk)�Z2[K��R��D���%z�4h-ѫ%z�䬖�բ��E��7V=[K�F^Bo�[����Z
���֢�E^o�XKkIc-Z_�i{��ٺ���f{��Z�XKע��E^���Ս<Gww9�yU���%zu��sڢWK�R���K|݈7�9Z�k��Zڸ�7r��Y@k)�Z2[���9{r�����4��ٵ�q-�_��.�r=j�Z�WK�j)�Z�����Z���%*������%��������kIc-9�%g��u�7� g��l-9��.k�^-ZKki�Z�,����^-�_�X�ۺ����R��d��"�E7⋼.d�_��>�Kv-ɮ%ٵhP|���p��ER��T�F�˻���E�㋜��t6���)h�Zڸ���:�����"�� Kv#?4H���ki�ZgK�l��Z�C�lɒ-��%8��}-5^KJl�-j_���忖���Zڸ��ג�Z
���ג�Zڸ��/�qD���.��tv-1�E%�\�:������k�-�[K�k�-a�Eq�\�"aKg׍<G��f�%��������$�n�셽���%�u#NHKآq�E��ږ[�^K�k�l-�[K�k��Zz��d�ҳ�ĸ�R�9�K�f�9�;��ג�Z�^+�d���֒ٺ��w���Z�=���'��l-:o�.��F?��z2[��*T\�dWHv�dWX�x#'��k!��=�Wh��V(�
i���
ѫ���ó�B�*�Y��c�`B+��n�Ʋ
�C+�^�CVh��U�Y�PU��
	�y���B�*��B�VU�PU��
9�Ѝ�,��Ս^�*��n�岲�0�B*,/MUa-a�F�Z�y%x�	���
A��z
�Ta�`B����\|�Q!��L�]*�B�)TI�*�yڮ!A��.�Q�]*D�B�SX%RO!�RO!�RO�xUR�*l��G���X�?��TB��K���
�P!J�n�㈞���PUU�PUU�PU(�
���
T�p*d�B6*d�B�FN����
T!A�Pa�⍜�YU蠺�SuTKj�B�*$�B�*�R�PUh�
9��
MU!AT!u#�r����Uh�
MU��*�R�PUU�PՍ޵���,��T�K�����
�Q!Tv#�ި���pm��
KC+lPC�TX�2[!�
�n�XnҪ�B�T�
�C�+,B��Gt��
)��)��
�CUHv�݈7�1���Vn�b���W(����rm����	a��1�n�X���.�Z!��X!��X!z��n���7�B֍�C��tզ��>�Pq�R�]i�Q!��B\*ĥBSU�K��T�K��y�5U��S/��R�
C�)�Bx)Ē�*��T
�S!�
�B�T(����p��8��I��� ;C6�FN��aT7��C�lT�F�lT��
٨��0�n�9�3���p0�R�킡�*tP��S�8�<S(�
��.���SXKv��q
T!�t#���p��e�BSUh�
	���
ᥐA
��J�B�S����B�(t=����J��>�sDI��T
��K
%Q!�z�Bx)��Bx�F�U+�"N7��2E�B�)D�BU�3�<S�tQH�(Q��(Q��(Q���y��j����pc=n��D!J��BUH��#����Z�%
Q�%��KԗXC�(D�Bn(�Bn(tP���.
�T�p*�®��
�Q�$*D�n�\�����Ѝ�N	�DPH��OX��J�
��P�R<!�";!�*�B>�F^/�D;�ʦ����B�'{Bd'DvBd'�s�ʾ��R<��)l��M!�R<!��9�y)DvBd'DvBSH���#���5$�V�2��	��9U�4�M��){B�'{Bd'4/����i���f)�K����I�H)@�4)@�4��F�!n)S�25)@��R�&ejn�Ty�KuF7�<��MJ���I�`R�&� ��M�AJ��R�&� ��M�AJɛ��I�E��(�lR�&�lR�&u��M�Ԥ��TT�4)@����&��\�Z�R+Qj%Ja��ؚR+Q��|N�礢�ٹ��gK��R�Q�$�R<)��";��(5�:��IuF)�s#��f��=�)�K=H�)��K�G)$��˥DP
��`O�3J)�Tg��RwQ
���M�ؖ6������I��Tg��9)��V��ң�p��R�Q��:���IuF)��";)��";)��";)�s#'�/5��(���N.ףOJ��9��Q>'�ȱ�k�K�EiG\J񤆣Tg�R<)ys#�P�Q�Ƥ%n��(h�^���Iј�I9��7�v���j�6(�OKMB�I(5	�&��$��,)�r#g�\v%eWRv%��8K*�яIx%��?l�ȩ����]I�n�X�&)o��&)o�Z�R+QJ�܈K��(���J
��pI*J�.I�B)I��$�\(���ɍ�^>*ʛ����7�ʅR*%��TJ�J����s#g�zAI�?�r9{w+A�T��+�#(�Jq��.Q�?)Β
�R�%u��n)�V�݈�j�[�J}C)�j�R&�`R&�^RGP�J�@)��R�O
Ф�LJˤB��I�T�25��'ejR�&ej����I����IA)@�4)�ֳ��?t!KˤڠT�.�(�^R!P*Jј��
�R��FN,S�25�#(u�%n)@�47r,�B��I��IU?)�.)���S�eiiYZj�I�<iYZJ��.��œ�,�e'�<KA�T��Gt�����ʍ8��JJ���I
���I���7Ie97��[p�*uR%EPR%EPR�NZ��R))���rRYN
���JJ����@�֠�pIJ�����-mFK��,-EPR�$�M���f�"(��&�MR�$�MRuMZ��֠��Iʛ܈�[��R))��"(7r�eʛ܈K(��v���st![��"(iOYʛ��I�I�AIK�R*%m K�ROMʮ��Jʮ��Ixg����SN�����'hR3N�Ԥ�h7�z�Ќ��qR'�TK��ƹ��{����I�����c�٤f�yDo�77r>�0NZ��6���ك���N*޹�'�/ؓR<)���K��N*޹����#œ�xRO��IY�����aZ�⹑c�X�x'�ύ�']<��'%�R"(5��ƞ9���7��'mlK۶��m�������l����g��ْJ7r,����C� [Ri�ض����Ҷ��F��ٶ�m��-p�����ϖ��*u�mf[ζ�l��l���R�F~s��`�칑���jp���y�Ev�Eb[dg��l+¶��-���l��mEؖ�ٚq�f�-��^���z�
n�6�-�r#���qK���o��˖p�.[�z�
n���-��Yn���}#������l7[���S�h��̖��zj�h��٢1[4f��lј��f+��
n��̖�٢1[�͖���2[Zf��l�5[f��l�5[f�l��9	��R�-���^�R�m�׍��Yf��lm6[4f�l7[f��٢17�Dcn�U�f�5�l���R�-fs#f/y�ej��^[O͖��h����@�m��Ji��_[O��S���l=5;\Ȳ>[�����������V���l7[��F��YHhKm�-���n�� $�m �jpn�$�Yf�S���lQ��g�m�8[���f���lm6[Hh	m!�muٖ��l��ж�l+��
n�����fKmQ���f�m=5[�h�mQ�9	~0����Yu��BB[Hh+��A[)��zj��жHl����ٻצ+ͦ���f��l�-�e}��ϖ�ق=[�͍�Ђ=7r.Q�8[�g��l����f�l���`϶�k�������";7�]VR<[�g��5�l)�-�s#'�U���x�f�-��Ev���m���y�e}�Λ-�s#���]"h���jp�Λ-t#f/��e}nļ{���y�Ev���-���ln�ik�ٖlm�4�ޭ��f��l�4[��V7���l)�9�F�g��l���϶��F~>�Z�%���][Hhk��BB�v��g���?[u͖���gmY���f��l�-�e}�n��[fKm��-����l��-�����Z[���|�Cף�Y[��F��x\�Ji�R���f�m���nf[f����DЖ�Ji�eV["h����c��'ų��l��T[�g��l��m'��ق=[��V$�{�n�yD�`��ٖYm���[fk��Pm{������VKma�m����25[�f��l�--���4[�f�li�--���li�-���^����@���Ji�h�VJ�5�l{�� ��٢17rx��q�)��VKm��� ����2[u͍��KT�e+��r0[fk����wm+�٢17r�6Wm��m����4[�fk��4�2��,g+�ْ7[Y����8[gK���s����n"���l� ���4�b�-S�ej�L͖�)��Q�djn�w^%fS
�J�O�Ԕ��yDn0%�s#O�̍��sJ�PI�����1��xJd�Dvn�is�)���)D���T�DP�*�B�\�l�*k�J�P�����s#�����r�yB�:JR�,�*�^*ᥒT*EE7r^<��M_%�TZ�J��F�y��JTRO%�T?Q� T	B� ԍޛ�lT�F������$�J+Qi%��;�U�.*�E���l ��׋����*i���*D%�U��J���+ѫ9/��B��*ѫRAT��
�9U�JΪ�+ѫ�*��J��+��*i��]TZ%�UZ%�UZe�X	h��*����*���ٺ��� �U2[%�U�n�}X>Hv�dWIv�:��*��*����*	���*˿J\�,�*k�J\�d�J6�l�*٨����û�d�J�l�*A��*��g*y��g*ᥒT*���Jt#?�W��RTT����9{�W�n��>�j8*uF%�TZ�J+Q��UbI%�T�n��]i�Jਬ�*uF7bxGe;W�3��^*�H%�T�L%�T�J,�F�>$�TJ�J,�ĒJ�QI*��ٻ	/��^*���d�4����pt��{B�e�o��L%�T�L%�T�J�Ψt��RTT���ޭyD�GuF%�T�L%�T��J,�d�J�PY�UbI%�T��J�Ѝ��Qэ��*��v�9/W��R)���ˇ@I�RAT�K%�T�K���$�J!PI��Y%]T�E%JTrC%7t#�rYY�U��J!P���G�*�?%$T��\V6W�❒��KO)�)���*񟲀���DPI�DPY@UBB%$T�?%�Sz}�����))��⹑��,Wn��ħ4��O)�)���Z�{J��{n�X>lI�|Ni�)1�ҲSZv�:���)����)]<%�S�87���l����~*��R�SJ|J>��sJ>�����ru�z�9{w%>�ħ�*%>%�S{J��{n�i�#u#���$�J���J��T��DP�#U�~J�O����R�ק$�J�ύ<!��SBB7�>����P��)U?7��ZSUG����J��t���rm���Ѝ�'>��ҟS�De�UI�J�*ˬJ���J���*��R�S�?%�S�>%�S�r���)Y�R�S�qJ3N		��P		�-X%$TA%TA%�SV^�f��)[�J���xJ���x�ʫ��))��)[�J�N��|N)�)e9��,�*58%�s#��_�xJ>�����#ys��m6G��H�����9�8G�H�ɛyD��ьs�l�����B>vx�#@s#�K�H�{�n�X�G�Α�9B/�ޭ#s�`�̱��h�9�2�v��������#Ssdj��̑�9�2GZ�H���NO�;���shn���i�#sDc��C��9�s�@7r^.Q��#�r$\����#������v!��9�#s�`��\������#�r�^����Jt#O���.:���Lͱ������+�r�9J��ң#fs#��ږ�9�1�#fs��G��#ysdj�L͍8�r�K�1�#fsdj�L͑�94GZ��˿��̑�9���#�������:�����9���),7��;��9J�n�����H7r��;�9G>�Fѭ\��H�)�c�׍�8���H�=HGұ"��A:�>G����܈I�7JGH�H��c)ٱ��F�M!xw?�EG���JG���̎j�#7t#��_Ɏ��:BBGH�F����HGG"�h8:�������yq\�����c3�%������cY�8:�EG���kЎ������fv���ϱ���.:BB7�B�+Mn�،v#'ᓻ���9Z��gG+ё��GtG:BB7r����\H��A:rC7�J���O;GG��(P:
��eiG��JG����n��rm� ݈#ڟvt*JG,�%��#�t#��)pt���ϱ���@v���I�D冎��#7tl ;AG"�HEEGQѱ��(*:�EG��H�9{��.:����#ptKɎV����h%:bIG+�K:2HG�F\�9�k���3����I��2m ;�PG�BmIG6�hK:ڒ�l�уt#g�OԂPG��F��6���H=�#�tt�D7r�>��8�ȱ|^-�W���ٻ��e%u#��:z����:J���gG��HP�GG���]tt݈�q|�<�EEG��XJv,%;���
�#u����q:Z���ӱ�� :ROG+ѱ��F�e���HPΎՑ�:��g�6�#u#���O��q:��mfG��8y�#�t䙎:�#�t$������3�vOk�4=H7r>�J=��#�$*u�� ԑz:RO�γ#ul3;j���#�t(�#�t䙎<ӱ"��3y�#�t䙎<�Q�tD����Q�t,;㖩-�Kq�#u�;�QG�8�#�t#�w=�8y�#�t�����^:6}I����X�u����]GR�H*��#�t#��w���I�h:bI�Z��\�FN��@ᥣ��F�zTTt䙎<�^:���<S�3�<S+j�qj�B-���L-���K��%�ZR�m�jU?-�t#�����k��L-���L-�Ԫ~n��᡹� Tk�i���zj�qj�Z�-%k�^��c��[,�ŒZ,�e�n�cx/�U���ҍ<!��V�s#ƒgjy��gjy�V��J|n�TycmU?-�t#���9��ݲ���j������Zx�5��ȋ�ڶe�����k-���L-���K-��bI-���Z��Z��n�i�j��n��Ǐg�8j��8j�@�קe�Z����(э�e���-Kk�V�s#���%jQ�%j��Z��E���c��-�9;�Z֧�崬O����ύ<�;��O���eimYZ���ei-���hZ���P۟v#/�{�(Q�݈ᅄZ"�FL"�m��sڂ���i����i��9/_��,8k�@-��
�Z��u����ͬ��6��ͬ5	��I�����P	��h�\��n�}B�j��Zn��Z�P���P[��*�Z����Z�P��P[�֢D-JԖ��(Q�.j�1	D7bx[�Z,�F�V�����Zx�u��R/��R۲�bI���e�Z���:�VgԶ���R+*j�Kj��Aj[�Z��E�Z��%�n�$|��J������v���V��j��Z��mYk�D�����Z"��TkuF-7�rCmZk%j�D-$Ԗ����VT����V��7�2H-���$�ܷe�ZwQ� �R� ��Kj��Kj���R�%�^O��ûIK*��R۲�J�ZR�U��#����p��-�\��K�s��I�3��R۲�|�FQ�R�3�N���홧�<�{��S�8���s���e�Z���Z���=����`������3��O�j٨���Z�S���Rm�[[��J�Z\�ťZI�S�y	���ݽ���ZΪ�Z�T�Y����Ay��:�ZyUKc���܈R^՚�Z��_�F��p��Z�U�l�֫���m�kɮ��MySЍպ�ZV[A׊�Z�#�<!����l�}rW�ղd�A�e�چ�k��V�ղd-Kֲd�.���V�V^�ʫZSUk�jMU-�բWm�\�^��r�]����FN�'w��z�!qUm�{���L�>�Kc�w]#��{�4V�Y��S#�wu(�z���ǽ��2��Z�}�|!�jѫ�jѫ���&^ף�VKc�4V�]�Z-�u#&!��ʫZf�e��:����5U�W�q�W�q��u7r�ma��ja�V^��_m�]����w7��x����:��ήe�Z��a�xY˒�֫/k��z�g-q��e-%�*�Z�U���yy��j�UmQ][T׶ҵ�XK��H؍�Nbl���[�F$lD��r����Fpl�^����k�F��F���X.7�e#^6�ec��X.7�ƾ�/uYc��hК,�Qq5ʫF�k4U���	����mla��ɮ9/�kGՍ^�k��F�k��n�$���	)���������1��1��g5b\��j,q}V��j�Y���yD�kG�k�Y���{��#�;�_���F��u�F-�X�6"a#6V���B���􈄍H؈���p#%v#/;�<�k[Jl��;�F�ld�Fy�h���A5�c#%6Rb��j�FS�Ȓ�,�Ȓ�,�X�6z�Fo�؟6�e#K6�d�Jj��F$lD�F$l��F��{���1����Pc����6�F�k;�2���mĸn��3�楑�ɮ�캑���7Cɮ��1��i��	�����c�:��F�j��F�jll��9�kH?��Y�2���m��F�j�g�K�yi4/���H=���X�6ROcc�H=���h^��F�i4/��y�`(��������ic3�(=�yB>�	�5h��hlF��K��Qg4�Fxi��:�q�q���m���#���n�]�z�Fxi��n��SGx�F��Sz4���Ӎ�hU#����3�-k#�4"Nc�ڈ8��ӈ8��ѩ4�Lcۈ8�<���6"N#�4
�FRi$�F��/��ٻ��,��KmI7�]�bI����F[��j������R�t#>mI7�GQ�%����J#J4�D#J4�D#74rCc�܈���Q�t#'�B�A����nd�F?ӈ%�ʦQ�4�r��n$�Fi�8�t#J4�D#4��F"h�F�g,��K7b��]��D{n�X>�j^Y��)�Ѽ4�8cw��2��Ϲ�SuY�l�M#�3�9��i�sF>g�qF�f�lF�fT6�����ȩ�`dj�ڸ��9�Qg4��ƶ���{/S3�F�f�`�.���9��xmt���]44��hh�^��i�9�__9��emDcF+�H���+�C`�%��mh�����6b6#f34���Fч@1�iwuF#-3�F�fhFZf�� ͍�� �Xw#'�;�L��Ԍj�Q�4�7#f3b6#3r0#�2.#�2�,�i$\F5���6B/3>J������6.#�r#��fc�Ȯ�%n3ns.�i�^F5�������������F��7Ci���јA�t���������!���_�����I���_�$�>���I�}x�6ro
��^���/���^����^���j���]�/r���/r�o
/���{Sx����aV����"��w�����~�c�]�/r��?�������_�	�}x������>��I@޼���Լ�K�S�F��ϵ@�"�r!��_���_��.d0�9����E���y�G�����A���}�E�U@�"g��a�E���"�хS�"�ѵM�ۋ<����9	� �������\�"�w!�ټ��]ې7/r.w,N/��s^ļ�s^�Tq=������I�@�܋<mo�^�9z7�\^U� {^�},�o�EN�'��^����b�"��g �;�7�Q/��)�z��pmcqz�Gt!#czx�ڵ��"N�z�1/�����R �y�6W�γ9/���8/�kB3ڋ���U��^��R��"����"���?�ȩ��A޼ȩ�[���#���3z�G�{�s#�W�/9������8/b,`���	y�".!��9����^��!��^�]
�R���"/��d�E��GE����Q8�/x�����{s��y�W¥ -s#��̋<G�B���x�nt���#�+�O|t��?�B/b^`67r�ټ�٣z��.+0�yD�Ӷ?� z��J��y���r�mW���?y�|@��s#�Eb/rx߭�{�����"��c�ˋ��[{^��t0���#�`（�y�	��n��y���E���F�4�;/r,�a�`^�X.>���q����yD7A��"����y�����E^	�1Ac^似�Ƽ�I�pJ�ً�����Լ�Ὓ�ټ��𞶿�`칑w \</��p�m����ʵy�"� ͋�=L͋��T���?����E\��y%\��]΋<�K��aj^����y���#,�͋��n�hp^�$\ihp^�$\|4�����]i4���s�_2�[9ei��=vx�)K{���O��y����9�%��I�>�ы�}�E�Xҋ8G�>7�n��"����"'ᯝ�^���6��"�����^�콛P��"��� ��"����n�r8z���Ɗ������r�Tz��'wAO��n�`I/b� G/b��E7r�B���:�!���C>�qu��y�û`�����~!�^��AYڋ<��јq����&=n�������~A�^���A/�J���x^�9�����E��[�����"/��"�E΋]�������Ź��s���>!�O"�Ì��C��"��r��n��~A�D�'���y.'���		}�r^��O|�s^�G�r��T{�׋���c��(K{я?��y��P�܈����$�>�;/�1�W���ß�"������|�>���'��I�|�s^ą�я�9Ǐ��ß�"������(K{�G���F|��>Z�^ćFڋ��.>�:/r��۟DЇe�E���c��(^{��rm#�y�Gd+���ó�BB.�y�<m�E�t�'$�		}{^��<ZBBz�9��]"���{>)�1�`�'���܈�K�|�����*���|�x^��ݷq����� �y�'�&��),~۾�c��Evn�X.d)�O�����x>
�^��q�.���χ��E~n�8�^�i�&�!z�'�#�'J�!z�û���n�T}rG�"���э�q�K�Xn��ږT�Ē�V�X.d
�^��A.�z^2�o/rx7||C/����G�ۋ��w A�O��z���n��)�F}��^���MQы~�WN��ty�ы~����3�<Ӈ��9�C��Ћ8�t����b{�F�*]l/�z�K}�R�l7�1�ы<m�m���z�y%\��X��9��5ҋ����E^�m�HO��$|���P#��k�5j�y�.dlI/r^.wɮ�^����>�{}�^�cx�ѭ\����$�>:����EL���1Uɮ���1/J/r��8�^ĕ�6�	_��KT����(q{�c��b8�����UK=ۋ<�K�ы~��Su=���"��J��o��]�_���'���}����+ႡR�ELUf�Ã�"��ׇ�E\	ɮO����P#�ȷ_<H/r,�L��wы��;���'���Y}BU�P�'T�	U�����*g��Y}T���'�	B}RO���W��r�kH6꓍�d�>�D/b��Pd/b,�n�9�DE/r^>P��"���������]�"Oȕv��D�>9�O�ꓳ�p��#��^}�WңyڮZ��O��Cg�"/����^���D�>G/�[�s�q�8}ԍ����-���qUE�>4K/�1<�(���S�"��Q��9��Q����=I>Zn�k��BB��Ї�F~�%�>ʿ^�c,?���D:�y�nM�>���G�׋�Mwы�Ю��!Pn��]�"��o�E\�q�$�"��[/r,�&��On�C.�"�r;��0	����;��>!��Ћ�8\ih�^��+�X/r��4�B���#�Ì�h�^�wY��|�=��9�F�g	�,��E�Ջ���xn�w�K��R���,��%-�Dc�h��Yr0K��R��h�z�ߏcQ-��L�x����{�h�̒�Yr0K3Β�Y�r���%���,e97����dj�L��Y�q� ��Y�2Kf�#�"�(���,��9	6�Eiԋ��|l'K�e)�Y
n��˒]Y�l�8˒]Y�+K�͒7Y�&K�dI,鏥�e�z��y�%���E^	���ǒ�X�_��%#�B��%�������^�cI,鏥�e	�,�%�D=���eigY�K�c)lY�Kaˢ��E^hW�@Ȣ��E��oi������C�K��Y�V�yڮG!�E�Ӌ��0K���XBK��F?��pՆ�V�c�z܈I�u,u3�j�yD� TK��s�!�EN�W�ECԋ���V�c�Y�K���<m�9!�E�ԋ��KT�c	q,!�%�q�U��1\�
nn��>c*�Y�d����-s#O�e%���3���%?��'�O/�%#n�$��F��Ēy���G�!0]
h��Í��O|bKb�A,��y%���_ra�%�d���pXK�aI3,i�%��D}M/�1����J��-��,��^�Xt?���8,�%����R]�T�,��%Ͱ�~��+�
�9	�&1�%�huz�軕��R]��6�%�dn�G���fIF,Ɉ�]|2K��Rp���4�]Xzj�����fQ��"�>=JF,�^ļ$#n�9JF,��%���pz稁f�),��^�]|T8��?�����hOz��r	8,i�%Ͱ��֘%Ͱ�K/r^.��O��}�sx~'_41���X��K�\��7�U�,1K2b�<܈?��я���%����������9	N/EO/r^>�
^,)���f�T,��%R��ͬ���ÒyX2K�ai�YbKb�A,1��HfIF,�27rxף"��"�F���OE��X"�e*�Y*b��Ē�X�K~b��Y*b��ō8!E2K�b�O,�/K�˒�XRKE�R�d1�>��fizY�^�Ǣ����;{t�:�>�E�Ս��w �%#�B-X�=���z,!���eizY�^�\Ǣ��E^/�(5U/����Y���Y�_����(�zS��XZcn�šG�F�,*�YTK�ȱ�����r�,E2KFdQ-��c����B�֘E�ԋ�_}B�@ȢG�F>�J,�E�ԍ\��zT$��,E2KFd�@=�Gذ�)BB�ˍ��vX�_B�K����P�b#!6b#7���BaKX�t#�g������B;Kț��I���&�m.lu
[�BK�]	y�.	%+!or#'��
y���)�KB�$$IBl$�������B��FN�_j�s�~<��Z�1/.a9S�p	q�P�r#�&B/!�.7�Z[�B�K�p	i���	9�yD~����]	%+!�zWn��C�%lb��'��֨�2!-s#��2�X
���x��(7r.>ј�	ј�	])a	RЄ M�O	�)a	RHބ�M�ԄLMX�JVB�&������	�*a/RHބLM(Y	1��	1��	�+!y�77�<��0N(l	��n��q�FN��Cd�F~}yh�,��%�xBˍ<!o�Wݐ�	Y���	��BaK����O����ύ8m���	�,!�R<!�R<��%{B�K�u	�.�`4��DP��	;�B�'{B���������	�,��%�Bd'DvBd'������	��9U�ܭ�
�-���F�e%��=!�s#fo�T�b	U,�w%���b��G*$�B"(T��O(3	)��o�MB����{%���_rY��m*�B�I�6A!A!A��F��PH(�n�9������P��[�W��hQ�ЂrC��$�
k�B�IH��U!]�E!J�?a�UH�5U!��T�~�
��n�p���(Q�����+��B�J�]Y�w�F~h�MĒb{�K
颰>+����Q��Q�b	U,7�z��$�BK�b	�лr��{B��B�)t��XR�p	.!�Vq�ȱ|�^
�-a�V�8�*�q
�,7����%��BaK(l	�P�r#g�������g٨��
}0��%ĥB�KB��SH=��SH=�>��
1a}Vh�	}0�&,�
A��
�17r�.wq�P$T7rx��UHP�Uػ�n��T�F�lT���P!�P!�t#����S�3��\���?t����S�3�<SX���W�)��
�B*�n�c|���F�P$�R7rxףn��
u3!�dBkLB� T�8��S�3݈�Ƅ�S(�	��B�LB��X!�t#�r=�\u#�r=
/E��
/���^+��Y��ҍ���.>=57rns�J���F^	�}E�BOMH=��U!��kB�)D�BuM�8��ӍK)͍k|Еz�'$�"N!�
nB�)tބ�Ya}VؕRO!�RO!�"N!�bIa�U�/�2H!p�kB�F�岒A
�4!�t#����&$�n�$\i�K��&�B�)Tׄ<S
/��^J���A����N���f�vR��T)���Ji�T�6�2H)���H���XN���Tps#?!���G*�J{�RR)%�n��y3L{�R��F��6�"N)�"N7���R�)��S�8��R7r,�^J颴4*?��tQJ�(Q��DPZ���?)듲>)�
nҾ�Tp��3�DP�ĔBB7��n�rCi9SJ��K)�Ai�R
	��I)�A)�ZvR�N��IQ�y�y�K��yB?�)]�BB)���sR�'{RYN�줲�T��";)��jpn�\V�9)���97��\�R<)œ�7)y��rR'�qR�N�٤��Ԍ�25)@��rR�&���F)�r0)��B/��&�`R&-.Jј����L
���Kj���}�F���gIٕ�]Iٕ�]Iٕ�S��e�����J*�IE2)�r#'�R�]Ik�RP%EP2\
�Ꚕ]Iٕ�]IA�AI�47�z���*�~ɵ٤6�� (-J	�Tp�.)�.7r�cv*������a�OJ��8K��Iٕ�]Iٕ�]IK}�R��f��+��&�KR�$%IR��F���"�%iyN
�����O�F��+M��F��Ꚕ7I=5)���f�֝�b'��I��yD~^Ky��7I��S��$)I�2")#��)ꑺeR�#E=R�LJ�\G�u�;�n&�:�֝����p���'eDRF$eDn�\�!)��lR $Uפ�H꩹(�B)đB��&�ҤxF�g�xƍ�#đB)đ)eq#�ЭIM�O��D�O��D�Oܝ��]C�`R~"�'R~"�'RX"ɤ�;7r^�V�D
K܈s���F|���&�ͤHE��IE2)?��_R"m�I�tR�KJF���vY�����DZ��Zcn�	�[IF�>���HɈ��b)q#'���H�17r�Z���HɈT��`RX"m�I����H��yB.Q�2)x��dR�"�,R�LJY�HE*�IE2�"&պ��}	p,W�dDJF����Β27��%#RK
K��DZ��)q#Oȕ�.+Ɉ��H}0�&�%RLJF���HɈ�������>7��'R~"�'R~"-J�2)R��)?�*bR~"�Jk�R�LJY�HE����T�HEZ#�Zcn�X�m�1)��Zc�f��F(���#���xS�l(ɤ\G�,��@��F��r�Y(�8R�LJl��C9�m��n�Xn�r���F'���lQ�-ı�8�Ƕ�hqlu3[�c�ٺe��V7��:�\��-��7�B�ƣm��V7��?���-�q#g�&��8��H7r���۪���f�l�-��u�l�-���?�6�m{���
nn�cxϑ��b#�B��g����%[���y�u�l�7[e+�ٖ3m�7[Pe���#��o7[��Vp�mu�
nn�9z��i���,7�)�״%\�����f�״?��6�-���R����ko��.dq���fK���stm���eWn�X��ɖ]ٲ+���?gK�l	��Rg���V�?g����%��f��l����̍�� �^.de9[Y������'��,g�l�8�N�-����lɛ-S�ejn��<�o1��g��ْ7[�fk��4[)͍<��]͖��25[��F��w =5[O͍���])͖���9[>g�lۦ�0��Ss#�w�+��h�0��5�lۦn�c,���@��xn�Gk���_ۦ���VJ���l����R�j�y%|&��zj�DЖ⹑û�5�l������p�YS����Aۚ���fKm�5��-7�冶�Ѝ��Λ-J�-���E[nh���#��冶-X7����U+pt#>G-;�b�-����]Y7�1�����X�8�jp�(�V���n�$\�cm�87rx7V��-pt#Oۅ��f� m�m}�K�:o���-��m��V^m颭�f+��G�ʫ-p�����֌s#.�f�9	��X��y�Œ�X�K�bI[uͶ+ko�<Ӗg��ûj���Λ-�t#���.����f�8m�-�Œ�R���fmu3�b�-7���lQ��HfKm�17r.�rOK�Zc��Ѷkۂ�m�����y�\VbI[,i�%m�2�ޭ�[fۻ�噶<�V$��l�m��V$�E��<Ӷk�8m�����mWֶ+kBmA�-���lA�-���l�17��Ee��U\[\j�Km٨-��U�l1[E̖z��gm�1[E̶+kk���R[\j������E���������"�mW��-�u���I������*b�lԖ��*b���-�E��<����噶<�^��K[,i�%m���f�ْJ[����r#���a'ն�j�p�:\��m'Ս�mN�i�3my���e[S����RO�N�-ϴm��"N[�i�3my���F��e%��U���K�c�֘-.�ť������R[��}\�]ȂP�~�-��%����}@�}^U��-��bI[�˶�j� mM/[,ikzْJ[,�Fх,������V�%��ޕ-ųm�ڂ=[�g�b٪X��������j�-�e}�`O)l)�����*{�J��F/����Ƿ��~*ɛ�թ4��0NIޔ�O7r,އJ�JIޔF���)ɛ��)ɛyq�;J̦��+� MI˔hL���EO%�R�R��z)	��xf*])%�R�+%�R�*%�r�cq%>n�Q�UJP�U�r��])�,7��%�R:\J¥$\n�Gk�S�u)9���)M/�֥Ժ�Z������୩����B�)1��)����)�,7��M�$\J���YJ��dW�V��J)[��
��])ٕR�R�:�N%�R�,%�RR)%�R�_J*�lu*}0���Mʾ�RS"(7r,W�pI	��R�R�%���F^	o�	�u���yE*�/%�R�*e{RٞTR)���J*y���s�S"(%�R*bJ*�TĔ��A)17rx�_{�JP�U�^��])u37�]�v,�8ˍ<"�K�)=5%�R.����^J�lb*��J4�F~�:�en��q�V�S25%@S�2�?�hJ���en�T�O��ȋ������M�ٔ�͍<�� �7%yS�7eCT�ٔ�M	Д M	Д M��)����);�J̦�lJ�O)��;Sz�)ɛ�)ˬJ�OYfU�9%yS�7%yS�`�����Sz}J�O)�)ۦJ��l���){�J�$oJ��FNյ���dj����Sz}j�X����lJ�O�ٔ�M��)����)���)��J��djJ�O�#U25��hʆ��!�djn�]ib6%fs#�r��ԔLM�����v��7T�7%fSb6�\�,�*ɛ��)MB�I���#����ڠ��)�A%�S��J�Ѝ���	{�J"�F���P�#U��J"�$�J"�ʛ�V��4��DPI�DP������*��9��J̦��&����ɏᝪ+Md�DvJ��qJ̦�lJ̦���K%SS��J��4	���n��ʅ�r��$T�7%fSv,� ͍�^4%Sv,��s�{�6�F��gL1��)�����c��LI���Ki�)�?�꧄^J�OY�t#�����@)@S:������M�ٔ�M)*1���)�R�S25���	)*�@7r�V�.��K�6��]����é�N���N� ��ûj%oJ��F^/�����K��O	�0N	�0N�ԔLM� *1��)i�9���r�R.Tb6%fS�3��M�*ɛ��);�J�����^���Sz}J̦�lJ̦�lJ̦�lJ!PI��ȩ�K�ڠRT�5��N���Gtm�*��J�Pi*MB7�qD?׶(QYU��J�Pi*��:��T*��A*����Ē�A��Gt!�U���ұ!��u��A7�{�Gmб��c=ʅ�QG��Xu���#�tTDG��H=�ci��$tl�:�LG�Ѝ��xl�:ROG��Qt$����c�ӱ��F��z���^�#u�����Q�s�����c�ԑ�:�~n�$T���#Tu���P�Qt���P���s�����p��^���4������B�\�BUGm�Qt$����:�Q��#�ttˬ���^:6W�AG��(:RO7r�m�@�~�#.u�	�yڼ#��#Tu$����c�Ս��^[���Ց�:TG6��9�~���#u��ƞ#u4��=Gcϑ�:TG��Q�s�+�ʫ�e�B�#�tt���\|"N�ʫ9U� �Y<�٨���K%>G\�(�9J|�PՍ�����Ց�:rVG��U%>GcϱQ�HP%>ǒ�#.uĥ����:�P'x�=ROG��H=�>G�B��l��:vx٨#ud��lԑ�:�QǊ�#u������$t���ck؍޻�<�^:�K�>�#�tĒn��~�X���s����#pt��(ё:�)7t#�w����#�s#>!���z�#$t���DБ:邱5��%>'�~E��^�#]t�;GG���>7����EGc���s���#7t��]<�>�qD+�ё.:z}���Ѳsd}���q���-;G�΍�ŧR���e�H���=!70��#7t�����:BBG�Α�9*u��џs�s�|ΑϹ��r�����#�s�q�M_G>甋O�(�9b6�|��я?t^.�;G����܈�x�H��ĎEbG>����=G=�Q�s�;{n�T]�AGc���s�);J|�(�����]T��9�w��bG����:�n�yD�����#7tt��;G�Α.:�xnļ�n�$���Q�s#����n��H*�@G!б�h�9�L���#�ttAG�H=�AG�F�F\�F~\����j���#�tlF;
��B�#.u,K;
�����tlF;T�?r>4U	�#Auĥ�l��Jt�.;�L7��KG��Q���.AG����#���:2HG��K:��n�v��g����qX��q:"NG���3y����زv�A�#uT�U?G��^:v��9/�}��Q��X]v�.���:2H7��_9/w+�?GR�H*��#�td��t�Q�s���t��9�=G��F���|�=7��$�sl����ˢ`�Q.t�;�=Ǌ�#�sl;�>G���7td}���QAtl ;AǺ����%�n�w�VAt����ZQQ[J֖��tэ���<"/�m)Y	���j�H��%����n�%�Z֧e}ZQ� j)��ë{n�	��ZQQ[�նs�O�紘͍~��SejK�nĕ�iɛVT�25-S�25-S��Z���eZZ���V��J�25-S�257�RT�b6-f�b6���F�#������V�V.��z��N� jDm;W����8m;W��|΍<!��΍��Y��q�cl����i�Z�%oZQQ� jK�ZZ�U�ȱ\�*�Z�%oZ���j�D-y�b6-f���(fӊ��b�ƹ������]t#/��OwQ�.j���i���i�Z��EvZQ�Դ M�ƴ�X--Ӷ`� MK�܈��eZZ�EcZ�P+��Gt����LK˴�L[y�j�n��]i4-@�c�LM�Դ MK˴hL�ƴhL���L���Gt�i�@-�:�Z4�FN��Dے����Gt3��iK�Z�����%[��%on�i�����qZ!P�܈�qZ�U���Mk�ia���i�=m�Vk�i�ڮ��i�>�ק{�F���ia���F^	~jɛV��6j��Y-f�25m�V�����EU����N�j�_}Z�O+�i��F��⹑�w��i�?����xZ���xZ>��%[m�֍�8����O+j�?-���g_�>-�Ӫ~Z�O��iY���i���i��Zd�U��z�V�s#�w��i�<7rx�L%>���F?��'�B�j��i�;�x�{�ޭ����	�v��i�=�����ZcO[��{Z��F\{�ZcO� ��Q+�iQ�jY��w�{Z>��sn�cxOۍU���sڒ�9��V!P[��:�Z����������m�jU?-��z}Z֧�xZ��%oZ̦����M��i����iU?-S��Z�O�Դ�Y��� Mд�LK��q=
д&�9/tejZ�Pkj�AmWۻ�j�ZmPۨ�257�1��胮�MK޴�L�jј�iD-��.�����%[-��g�ƞ�+���j�;7r,�z���i����i%>-f�b6-fs#.� Mд�̍<G�49�V��{Z¥eWZv�eWZv�5���#���ħ���hL�ƴL[y�z}n�	����i�>�ק%oZ�O�ٴ�M�ٴ�M�ٴB���i�Z��ejn�i�jɛ��iA��%on���F���j%>7rx�9U?�קm�j���i)��i�<-�s#��S���x�"��i]<-��R<-�ӺxZ��EvZ>�%oZ=O����Fg�qFg�qF���0����Ip����3{Fgl3���%>��gDvn�X�#�s#?Z� ��g,8�F�g����ύ<!6��Ǫ����3A#4�X�#t#���:BB��gT��(���!���3A��gt�Ѝ�в>cu٨����-Բ3rCc��Xp6BB#$4Acuٍ���F=ύ�8<4�.���3A#4�y�R���l�Fnh����K�B��3BB#$4BB#�3���z�Q�3A#4�?#�3�?c��H�ƞ�l�9j����f�Q�s#N[cύ8G����3z}Ƃ�%Q�%%>#4�wn��{#��z��3�>#�3�>#�3�y�ۃ�f(�3�=#�s#g�#�����]iBB�xg�FH�FN��r˴�l,%���:#�3�?c٨�!�Ѳ3rC7��E�)�9U7V�ь3�>�g�F�g�F�g�˿F�g�U+�3R<#�3�8c�׍<G�c������_7r�ZY���)�џ3�=#�3�=�>����^#�3R<�Rg{�F�1{i���58�g�ٌ���~�ٌ������ru(�m6#y3�7#y3b6c֤�{ј��j�ٌ�W��f�`Ff�__m6#�2zjf��z[�Ff�^n��݇�Ҍ�U��f�Ԍ8ˈ��8�h�	�Q]3Jif�`�YF��	��p	���j$\F�e�YF�F�˽c�"%�2zjn��W$q��]4#�2�*#�2R)#�2R)��ވ�j��k:7r,W���Ȯ�Bi#O�'>-;�?g,��7��f�ٌ�����Q]3�1#�2zjFO��9�W.f�	�[�k�^����r!K����W,b�X.Q4��f$\F����n�z��Q73r0�Hf�YFvedWFPeԺ�������H��T�(�/#�2�_F��hz	��p	�g$r=*�yF3"�"�z��z���p�2�[f��1��el�ٕ'��˪]Vj]F�el�M/�����D.+	��!jt�����2"(��e�MF;�hg���J;�Fa������]y����h��Z��QD�0�XFeT��@Ȩby�~n���y��kļdDF���9"_���t�����p�U,c����@���4!��e�~��[�n���&2�^�V�y�Dn�^F�d�p��[�F��(��+�F��Ȉ�Q�22"��e���������?����#�Y��ߖ������߲�o�k�s^?�[?���{]�o�c~�c.�c.���c������t����c.������8F�8��q��q�Ώ���1��q��1�o=�7�q��y����c�c�c�ϲw~w~\��q���͏�̏��X���r�o�5�~���!$�͜�����d����cM?���c���$�o�c~��\~��� ��~��cM��o���Z��R�ُ�?�?�?������؏�f?Σ~�G��K��~���~���|?����0��~�������������~���cͬ�����f�o���֏��?��3��?������f��d�7�1��1�����׏5�~���c_]?�����G��7�1��q�{���1��~��>�?������'�{���u�~����\?����&��~���\?����׮����������_�{c�xf�{c����>?�y�x��?���=�{c����uu����(�BQ�H�Z�T*� ���AGP�fܜ��z��6��f���j����7���>]������_-�[��
q��[?*�Q!.�?*Ĳ���o�3�XV����w��X��ϻp�1>S��Ƹoķ�xnĲFN��	1��~j*_��^~�ǆ��x��<�1��1�q���5�xc�7�xc�7�i#k�퍱�ȯc�Q[5b@#��L�6�ą��������@^7��~`<�8�������@.50��R��@��2�6\�00��Ruπ�Ċ?�<l ���m V�\uπ��@����@-4��:{�|u�@<��˸�o7����O������~���v>Ǎ�uço�f7r�1�F���7�q�/��7���Z�F�tc���7r���_��7����ߍq#F��7z7|�Fv�?n�����g&|f"���g&bބ�Mķ	?��	?��߹=_���'|k"^N�Ɖ�p���>�D\���y�Dl���&��D���M��D�8�矈o?��k�u'|"��&�Ӊx91GL��D|����\t"��E'戉9b����Ń<���?�Q<�m��?�����������W��x�������� g}����_>��=�>����-��>����ۃ�� �>��|�A�>�������䅸����䂿-��B~���.��B]����_.���\�9|u!�]�m|z�b�B]�����?_ȕ�|!v/Ժ�|!�/��Zwa.Y�u旅�e��]���:`!?X��j���iaZ`򃅸�07-Կ��B<_�7�˯3�p2�v\#��l���:�� O�i��{�\�i�:s����e�p/��9��u��f'�s�	0;q��|\��9o�u�ۦ��s�sD����#���.(�m���5�� ?���:�m���9M�
�Bq������\%�3W	�Cq�}� ?���P�
�Bۆ랹J�
�BV(��i�P�&�C~(���m���9R�+�C���E`�g��*0_�G
�H)�U�9Rę#E`^˴_~�x� ��mx6�k�y-0����)s���9q�*�)�2E�}��3/	�LF)sN`�	�9�9'0��YGE��~��߄��o�<�m;�i�/>�)>�)�2X� ������I"�$|�Q�3�6��9�� ?��.(���H�B"N'�#��8�m���}� {`�"�E"ւ=
�GQ��������UȽ~~h�p������B<*���(��`���3`�LѶ��S���(��CV(
�~(
�U��|�Q���G`�����ه�G���F�i��H;�9�U#wl�أhĞ��G��o5�Q���-�h�V��Q��	�_���7X�h�(�M�)>����A8� �vj����6bT���Kب �|S4|���Aŀ�ԃ`�b�/�Km��l�d5lԶ����T�ۀoĲW`��{�����`�lT� x� /�lT��8רlT����88�O��
�R*j+�M1��9~	�)n������70O�)�-�� �7|�F|��[`�,Sܨ�n�7�����[7r��v÷n����7z7|�F]�*�Pō<\U��pU�*n�2pUq��C7|U��
pP1�3�h"w�qk��&z�`�lT���6�r։�o��/9�OO��	���:�c��_�Q*�A�D̛�y`�b"�/�T���	?��s�R6*�A��m��"��K0O�)&�+&� ��m;��A��z�`���|����/���|W�F�|kԈ`�lԶ���A6*���|�y���A�C�m��`��O?�c�P8� b#�� ����pF��3`��Q�=
�G�0��8�X�G���Q�)
0E�(��B�?��b!n�
pA.(� ł,Ĳ�q�'���B�Z�[�xb!��	�9��O�ŉ�X�G����m�w�`l�:}+�3�$X���`qz7	>'���u�e��I�9	>'��W�N��I0;	f'��O^g-�`{=y�1/�ۓ������#lO��I�9	>g�pg�J06	�&��$ؙ;���I�3	N&�3&8���N��I�3	v&��$8���N��Mp2	N&��$����N��Ip2	흄�ζ�^0���I�3	v&��$ؙ�`]�K�uIh�d���ۓ��I�3	N&��$����q�����_�>��W3N ��mx�3Hh�$8��3?�8�;��J� %��mÿ;�m�s��E�heb� w��|�M��ٶ����$�������A��$8�Ǔ�$J0;��#�S�`{O��I�%؞��PBW(���w�	��mxWgΟyֺۆ߃�'|�B	]�S���\P�Y$8�Ǔ�Jp<	>'��$4�?	͟��O�����x^�U�m�1���%��,�`��D	�(�S��J�CۆgC</�j�W�%��������`��ϡ]�m�b|�ϡ]���<R�=JpF	�(�%8�,�~!��3JpFو���G	ݣ��m�؀RB�(>�(>-������H	-�g����Q�3JpF	�(�r#/g�`��P�ʆo5��/�/�e�/�˔�eJ�G	�(�e�=�l���:J	V(��P�J�C	���R�3�6�b�@{��B�)��51�m�{F�
F)�����r��5��
)�#%x�����<R��@~:�o��Ѷ�^P��=Jh5%4�zKۆk�����d�RB�)�ߔ`�ZMyc� ߔ7�s���`��S�ȁ�A��بm;�ب��S���6<|lTB�)�<������࠶���Rۆwz�R	ͩ��T��J0T	�*o�_pUۆw�� V	�*�Z%��U���6��`�UB7*�U%��W�`�U��J0T9��TB7*����Q	ݨ�nԶ�cZR	�*'�4X���W�P%�m��!�N��D�ZR	�*'|z��A�D�ߔ��:O	�)�<%������t��:O	^*���t���)��b(8���~�6\��S�eJ�L������m��@�lT>���JpP	�)���>ЈڶsL�o��ݨ�nT>��|�������\U��JpUۆk �Bs*�9�ЗJ�K%���W��J�Pm�����%�����
�+�n%t�<׶�� �׶���R	,�}%��ra� ����>,�/�`��S	>,����Q	���ЃJ�<%8���S�-Kpd	�,��%�������zP	.-��m���~-��%���Z]gQВ*�Fm�q�έ�sݪ��ط��m����
L۶��y�p�[�-+�ef������Yof���΄�6�˙�x���TA7�����V�~*�W��
g���pu�>]�Ҷ�=��V`��:�w��O��
\Z�7۶����BG�����*�~vAϨ�gT`�
�ح�U`�
:E�s�
�V��*0Y&��dm�{�߂NQ���U�
�V��*hx�
�%ح�U`�
�V��*�#�p+�#��
�H>������m罀�*�W`�
LV��*��V�G*�#X�U`�
�8���j6���T8����T�
g�m�|�H^��<����R��*pP}��>R��Vl�����[`�
�G���{�m�*�7h!8��Yj��A8���R��*h+بU`�
zK��U��
g�����RAG��7X��T�V*h+U��Κ���T`�
|SAo���T��
g����fҶ������
:J��-���ymn����m����T�Q*�H}��R�[�F�jĞ�/༶�T��
<RA���#Uc܃=*�Gۆ�1���ў6��=�6\>-���o���
�H}��>R�y*�#8��T`�
�Q�=���YoM�T8׭p^[A��p�[���S`v�����W+�=ۆw _��PA��
X��ym��ST`����8���NQ�*�x��S�x
g���¹i���ԍ<|ζ�^�����6�3��Nἶ�S`v
�Gۦ��]��oļ9!���>R�*�Bۆ�El?T��
�PA[����
�PAo����S`{
lO�|�m�=#�Bo���T`�
\P��)�1W8;�� ��S�Q*�>ާ����
�H�p�\�*pA}��mx�#�m����?T��
ZMۆ{F-	Ψ��T�t�6�3�!pKF���T��
�RA�p޶��-��T`�
:O���
,Ӷ����8ۮ�<ά+�M���7t�
�S�e*�L��S�o*�OW�t*�L����T�t*0O�p޶ទ�@#��PՃ�	�Qݨk�m�?�/�
�Uጾ�U`�
LV��*�۷m�?�9`�
�VA���CU`�
�ֶ�o1���*�V���*`�
U��*0T�3��c5;��CU`�
�TA'k���[���W�Zm�����*�n��+��W`�
�VA���d����ֶ�9����*��W`�
�\}�U�
�U�|�U�
Z\��p~޶���G@���P�/�m���R^��A8�Z�}��W�
T����W_g��K5ب��T��j�}58����^ͮ��VCw��F54�[��A5��lT��j�Q�����5��}^����8+�qV^��j�R���ն���mx�g��`�z_�������j�V����j�s5x���V��jpP������jhb54��Xۆ�1��U5���Y֪�Z5��g�5X�m�s��pv\�L�����U��j��`�LV�LV��j�;���Vǹ���j�n5Χk0Y&��_5بm;�TC���Fm��^�u�y���C�m�;��t֪�k��V�N�*����8wn�p�4���U���6�� t���?J�L"��|���q����T�L�γ��8��A5����TCK��%�ВjhI5ب���Ҷ��0�q&\�[j��m�{��SC���Am��#���O^��K5x�mý ���jpUۆw�����FԶ�o{�Km�>����Јj�Vۆk F��jhIm�=|�����g�m�y/`�:Tv�q.^C���x5���6\�)άkpZ�v~ˆ�C_��s5���ׅ�Cs��x5ζ�6\>�q�]��j�\}���T����T��jhI5α�6��*X��U��j�[N��C�m��A���/�`��08�4��S���,XCsj�p/�/�9�Зj�K5��g�5ز�K�F5t�Z㼻�yw}���`��Q�q�]�Kkpi.���5x�G�Сjpdf�q�]Cs���54�YCs��9�`�g�5��Z�\�ƹx}���m�; �����Z�_k�F54��Of�qV^�#kpd}�Wo�%��k0cۆk�Wo�*���C#��v#^B7���5t��Qݨ3�8{���`�|X��6�-r`�A5���ρ��OO��DL[��
f���5���8+��}5���Yy��s5ح��`��U��j�V��q�^O��Ј�6�|u�6��y֪�Z5��k����Qۆ�Cn;�8S��_m���`�����1ZR-�����5��k0Y�s��RN��i5X���ZR���75�������RC#�q�^�=j���8��5��g�5�m�u��/��ZR��q�^�e���QC���
m�����P�j�C~��m�� +��~jpA���VS�j�25��+���\P�j�25���R�j�����LV��
m�u(X����z���zKV����`�Gާ��l�~��WpA.h�`��m;�1��0@g�pAg��B�� +4p����~zKzK�р� S4�h0h0�GL� S4�pAzKzK�� ?4��Bۆk�1y��[��������.h�p/�1�h0h0�-��O��Q`�������8�o�<��h�)`�t�8��h���g�`���أ�h@�i�3�t��8�~h��}x��g���6��3���>�L�LzKlπ�� ۳mx6�/4���m�5�||@Gi�콁����|y��g�pF��H�4أ�h�)8+o��w�h@�i@�i��`�`��t�X�.h@�i�l�~h@�i���h@�i�)8�n༻���Fi����w@#j@#j$�/�������ݨmó��5�PhI0T��Z|������t����o`�8�M�6j��`���@n�i���m�-pF��h5m���h�|��h�|�i�=`�أ���t�����~h�8�n�̺�c����������ծs�#��3�of��qJ9~�r��Q����;��g���ϸgx��|~�?w^tW�������_�����AG�ߌ_6�y�_��s�_��g�~p�RƏF����k�������|�l��\�������������1��[�~ǉ�����(�y�?
��/�_���q��W_����:�竦}����?�������)S����~>�o��%����<�{~�i�g��B�+�����<��X����7�Y?u��������a��_x��=��x�������_����ϡ �gװ�_+�7��7�}�����ߟ��{���D��:��=��|����?�[�����P^?��3�~�����2o����3�yK���3+��G��$0�s�����������h���-�ߞ�?3�c���w�^���ٗ�yKK��/��<g��x���럸�X�!����q��裲��*�qaV����]�F�G:�s�8?����?{!�-�r�a���s�����T׾߽�v'&�{�Se���R3���?��'���|g0L��}��]N�!��`��������� ��o�sٓ�Ը�L`?:����~~�w|����g�'�3��'�af�1�}@��-��\;L���oV"�ܡ�~�-]���`�y]��o/ƫ���X3ξ�L�I�9'��L_wB~~�w��%F����u��>�7!?k������ ��{��f����͕��@,�?ɡ��k0��X����2���e~C��(3��@��3�}<��s������Q���H�wW�9��'f�k��o��w�����~��A��gD�c8?\b,�y~�y�l;Q=o�=��������̓wv��{�s��]g�ȏ��'9�� ՘��DU��w�!��>�o��.��t����~ӭs�$����{���:o�J�-�q�k�����<#׮0��"H�W�IT����l�f#�{A:o����ό�]`s���z���3:j��,[��?��׈V�@�bާ��n>x��������:]���v�$�>C�X��@U����wU7�_ʫ�!Vc!�V���<
�k��7*�F8��3[۩�v��W+��_a�?3"�X�XZ�OF�1Ϸ�#�$S��g��e���2�O�?F��3��!�w�q��~r�-;]���9����s�<{%��<K���qK5ѦX������'+������A��V�P�d.���:�v��̬"QM�/�{8B7J����g_u���t�q�[�v{���.C�dk�u��wG9�k�s,�0�{�uV�������?�
~.�O�g���S�{D��h%�]8��|��y�B���_w��}"5z��;��o�'ݡ�=�>ob�>���T|k��ʓW�w�ك���
�]L�o)�-�SD����(-�F��gg|��=K��f��k�;1Ӣg���[�}�W����|���..`�m�1��;r�������P��@�e����4T#�yȇ-���t��~"'<gV�>�h������je$R)�@��(W_��Ә���^#��B��9��sK��񨟜Zj�=��pX.�_�\�@G�Af���W��5b��\EjIK�~�}:�����~�Ht'�9������VF�P����g7&/4��N)�h�\O����>�s��;��1���@>'�+U4]�H�i62�1�D".,;��ٌdb�$�֛��w���S�9��g��gZKVh�$L>�2�,�1�Q�}�9vu��ܺ���1Xm	4�v���������|祳X�ȷ�����~�fr`�zW60�,&�@������g��w�)ܞ�
1n��SX��0�#`ԍ�6�.sk��'+w��&�֘��j@څ*�g���$Ia��]�G��A��(_z0�S��0]�G6�ό砍F?$ ��(
�x!�'ڡmɘZ���%7�*���j<�/�Qo�����]7��z�Q�,�������v�~��>�'ѯ�Qa,����B�a'fx�hd8�ʕ<O��ta?V��@C#��G���Z݃8{�o{~��e���L��X�9�quѧ�B�7z���ꥯI�g�|����U����u�Z&����  -��׈Tsa�/���v��Z
��ϧ0J�q}!1[�f�z d�=�q\x�9��#� ͮX��ea�g�r�%<O5W�|�B5Z1���{H'�������G#���s��s�Pn��b�ꅑ��
u���ׅ�+P�U�c����<Y(1�M`�����X� A���޼�P9�9�V\XX"0?F~<��ЩU�t��5������e-,&~Բ?�8@>\ Q��[�nLk{�b�o0���Ȃ,\j�=��w���|��*[�"^�8v) ���{���� [�*������f��T^w]�����,��%xG&�L[��φ��-�ev������.����=����X��Z���}�5q@(_P�X;�C���S�]�<���Cc��*t��o�}��XE�������}=7�,e�;_AϿ�jYׅ�O�)�-�Su�¤�`�X]2��Y�X�ٞ��_���9d{1&�Y�?;�v�9��*�{7����Dhd������̢T�0�4F,���
�_�9+y>�9��Y�����$��RT({JGg�Fiy�5��%R����=xK`���~2�u��]Z��~
�9���qZY�ٞz�!^H�>mŅ��X��&���
�R,^X��P(��!�*4��*����f`��kԟ��G��|�
�c�E��Mw�꣝���<3��(b��G{�Q+ij|��&��K}o�E�D{�ƍ9�FD���.7u�
����XP�л�A���:ƶ�J4E�e`4ñ�+����0nLo�e�����?������?���tط-yN����-�Z~�q��p6�Y�s�|PZ����諶��yt��B�{71�����/�vR����F��Z/~���Z�������c�v��Xx6o_�m^tx�k��m� I��s�b"���w��q�9Dh��=E�C5����kN����
�a+�;sG5�$��R������_�2�P+~�Z�`V�R�֫y��DQ�ĺ�~I�}Ԟ��t:ϱSw��h������\�ٽ�JL�{gk�_I����h�|��)h�F�e�>yN��kbQ�J�=�P^�c���7�Y �'搝j��s�B��!�R����S��X<���夰Tt�)��R��Ⴏ����}����g�y[�j�*o8�N����F'j&��]v��Ҏ����xI=X�����w)��Ծ3�z�}�|Ē��U����R�#q'7\#���6���>\�Bߦ��O���F;�D��k�Kk�;=@[XHݵ�
�>s�w/�vL�X-�
@#�B����Q�.�-npK�������G�y���e�xq�!J�`��W/��� 8-X�@�c�Ϯ�>�%�(ׅt�2���l�����F}>{Md���z��z0 얁�.����0.l�~<$����~�5�F��}�ʓ�	^��~�w��tﭞ�T��#�<+�M�������4�%�n��ju̴�t�2�{'��bGLȯ:��.F0��~���>a��[�SjO-�%M��ٱu�û�9X`u`a��.��7�N�
��a�5h���W�ۓ�)Y$�`���V�5�I ��ίP��=U"%~�H���2�pq,7R����~\ b_#�>�ѻ�߷-�|�t
�	�u�Rr�&Q�����g��n��v����#xuOZYV���s��U:��[�QƂ��ۚ���j���ٸ��:����|�_J3�9����H޳/��C+�֋#��>�9�W����q@��N��`T� z� ��~���o�O7DE�¦�Wt�!�]r��˵[��S�����Ȫ��_��� ]x
�O�K�v�иnm�]7�z��3��o��wF�j I�=�hu�������E3|b������A��SF��D]뜓w�A!2P^͜7�´�>����s�c�l�A��,�~9�/����v
��&�u�ߵ(/�3���KmL�b�C�����o���D�vD�>Sl5ʝ���� ��Fh6b�o
С��9\ᛘa��W_����M
����<�#qI<?�>f`�^�x��[�����N]{��}��j����.��6Q�E
�S*�`���mhb���H�hKn�j7DV�$��۷�#?B�I��	ߜ�)=�R��O�hz%�P �4)���e$���e�LeV�;@ㅔto����?>\H�V�œ�󐱼�*�� =R�JI1̐
����@�dxT���G0�$VH���<7DZ^�����8kc8��ڼ�#/0ޏ�W�6`J#k�:44��,"�}��%E���;5º�#�$ص}	=�K��;0�́F���w��L����-�=}��x~�@�����C�`仏�q��J������)���=8y�a���O���[	��_f��W���9������/���B�;���.���zǻ�^�w����X�K���2�3��T�s�3��Sx��5�߄���B��8����{JO`�h*�+�¤:��U'��
�	]��Y��%(��ů%��%A�	%��xm�@R�5/���\�h��ȁZ&p�ѫ�eG�0N���vGmЀ�t�l��괦�x��wm�� еc�y������!�p��IHG��2;D�s��Y�h���Hx ���!h>T`u���G:�j/�#�N�'дf���г�y�G�po �o�+msu�j�R�Ė�	mɗ��:T���%�`^ZTJ�:�Q�{(�}�r�MfTRN@w�Ө?���j���n�?�����ǿ�����?����/��_����������������������˿����'������˿������������?������/�������Z�.� 