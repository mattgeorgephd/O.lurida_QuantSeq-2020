�      ��	��GQ.^�9g�̜�;3'{NrfI��dBd�da'��Eք�oI�%l�"VA@Q�E7TPq��׋�^��� ������O��>_���	��r歯��������~���1�����l��7u67_��0W��قm+w=��/|�m/8����n}�O=�/2��eݶ����~�l.�[���Y!��֗{��)����R�=�D�j}���?�|�]>����^>�*�3��M��n��7�z����߀�s��[��?��w֝L�
>�;�m�2G��z��w��n�sF�}E�pL�?!�g^�O�v��s��OVeA��+�s�Y�w	|�Z?�g���a���l)�	�'�|{X�'�҉�:�|v��B������|�H��_\?����|Tc�&߱�6�i����93����|ft��<�g�t6,:.Y��,���J�?3z�.�]o|�|�(�Om ��=�]���*�xN��	��x@��6�ꩽ�B��mׇ��	��R�o�ߧ���zx���Z>���m��R����t=�?Z�:��uxw~��k�s��鈻��XG?�ܦp��zO��Qy;�>�=����"��@+�j��v9�s};uL�ɛo(���������\ 7��]��V�?�ԇ��;���#��{���6�s�sO,���g?����[����L�E�9o�|���u|�7�+�?\�ia8����چ��y]�����U�/�K��o��>�_Y��Sߗ�>�?S>�+�����[�_��EmFr�uF��~w���W9�TaΟ	��r���~z�щ>���x���<"'EW��"��^��g�A9�b�ܜ�Gۑ=b�1��oZ/O;���?��s���)����L}~@�<���'�'�o����_�����yp�<��������T����>���g�en�g+��n��9p�r�M�m���vYy����PgL~6�w*�������6��_��x~9�c��:�S�������7��8N���bz,�o�=��i�m�c�:�[�/�=��ņ�G��aѼP>,$p���w��v�׎�Fp�ujg���6��r���ؿ��Ř��xI���9�?����ϛm�����-_G�þ���,���G��~����#��Ǹ��|��g�g��k̓���mW���˟?/�g���ٯ����E���z��\�'[G�#���v7�j���L'񧻼������B�s�M��� �q�}�D�Mp��K���}lݷmد��?���W�G�5^ʷ���%�� ]�_�0�����<ѼS}�b����6�s���?�mhE�k׊꫽�T���x��L�6Y,?����.��^�?��W�ύ�S��;�?K��Й�=��6-?�CQ�,.��Y�7ǘ����@��N�+���*���|s��������@��ǆ~>��E��½���7�+X�d��,���ȏ2�<j�2��-6�з�b�������N.��)<��k||8F��{�l���{�o*�9ِ�6�ofH�t��ߟ-��/��h�E���j#�p��K���Ǎ�9�~��볷�qK�0'�]�Ga\7[����O؞1=3�'�<B��/�կ�8s��%n	�tІ�I�뺌���Ϙ�/W�1/��Y?︿���.��1�3L'��l|O�ϓu����7�&�f�Ѻ�b�0£� �.���
�u0�%�O?�/�ò}<��}[��z���G����й�}ջ?���Ŭu���&�!��=l8.�+T������>�'��M��nYG+�H�}����q�fA��o������9��&����i�W���8X�?��;�7:�u��Z�I�2>=R�㳊����O��?�?�\)8?��,�_�;�Ƀ؝��*�?U>�o��F��7�瘃���>��t�� ���o�~�8/���.�+A�,ޮ����绬�?d=�grnT��"�����p��p����0>�_��G�u��������˽,����
}����%|`<��X�[�=��py������/>�W�g�8�'Yϟ�۴�H�N�p��:ߡ϶�8���n��������ubG�Pz4�j,~2K��~
p].�����.�n��Yw9�!���K	����G�[�g�d� �K���]a��>I�5�oZ��|����?˜���<�ɦǷu>fyJ��\O�#���M��6�G��R]n��d��y��;2;r�M��cl]G�>YxO__>�=�E�P���y�կ`����q���!<l7��:&RE�����������_�o�j�������]�x-��?��K�$���|�>�|�,���>�;�8.Z�z{�:_8?'�/ʟl�˸l>��rw�hA��������d�kt�'߻��}�c������]���6�@�x/~����R>o�uyR��3M���i�O2}������!�Y:���F�ˑ:���q?��R��ɧ�r^�}�D��4���x�W�9�ǃ�h�8�E�
�>X����u������W>?i}���Y<hW������ҹ�����J�ϗ�|,��U/�<�n���[e����љ釬�ί��w��G
�7�?�x�w�N�x�t^�T���(�P��u�������.p�2?�w��!o���hE������.���<�_C��u�ש��ߎ�q��=�wP����F����aن�Ԁ�t��\�u�7�_�p��x���W��S���㲘��D�h�~z�n�l�^����~��X��)����M�_���Ň��ou�n�a�sU}>`��W�g�3�u���p�Ϧ��y���i����#��͆�q��'��c~�5��'�{K�km�����s�����&����� �������/���ay�d#���g��F�iV?��|^,�4���'���"�����-t����o:��+�گI}�}a��k�O��?��҉�c�O8����潻��U�r���yE���
�p�w��脝��~�����s���w)?��{�s^�3�Ńg�{o�����ϊ3Dz#���ɛ��x\����ր~�������Y_d�W�3�3����>�G��:��|H�~���x�q'���|�rZ@��	���
�x�����1+$�o�_���Y\1��t�E��V��͋�<�6��ȭ��|7�o�>���1�7xV�]��l�/e8΅��Z�0<���y��������$^w������9�V�����{���Ef/4�Ɵ_g�|���Ԫ��������w�8�W������u���|~#���O2��Y�,F�x>tY'���������Ƶ2����ev6;d��y9V�ϭ��:�n�����o���t\8�����\oG���F����*�evoP_�w��
��y����6�+��fz2=щx��-�.��xXn����o~ن�ݺ�p���X�]J?A�����m(�(̇++��z���d�K�8��]6�_F���>'xP7�+���b�>+{�~K�?�=E��H����ߩ|f~��A����Xް7��%�e9|~�������	�g|V}��oW��O�*?3z6�w���q�y���C���D��{~�E�6ˋ���K��3�6�
��cv-[��d�y����q.�����?�[�OG��H}��l}�%�3��Wb�v��S�h1?�v}��	�~2��Kb��3F�Sh��b���OUް�|ޔ�G�����:��>�O���S�9e��k��U�������k#x���8}���ѽjj�J�:�e{�	����>��2|���p�a��ǀ�?���}1wci�9TR��O|ݧ�c?��L/����@�s��I����r�F>�돍د,�[�w�龏���s1l�8�H����<7�=����οǹ�U��������y��������w�=���(
��}��l�d���6�'Y��_�S�y��=޷��{x׬���,mtWY�=�Y|���X�G/�J}�s;?�)hW�ǯXb��s^T�d|�B�F|���rt �����4ޅ�������}�oz`#�^j<��(>l��i;ۦ��c�j�}پC���E�~�o;,>��W��֏��w�k���4�ß������q��$8�7��+��D� �q�Й�_p_#����z�z>����Q����s�\Tn�����켼���-��f�͘������|~T}�q�W�'�`9_!:�vѶ�ǣ�Mf��q	E���<�mk~�Ϳ�}⾎���փ�?�/��
{���Ⱥf��D9��}fA��z��C�s���u����r�X��o�C/����G#b��D��y�xm��������nr��w�~�ǁ^$t^i=�Z�y@�c��y_��=R����|�?���Y��:^-����nw^k���<�~�.g�b�'��%�~�WW��F�*��q�?���{6-?��s�ED��!�#B�\ ������_Gp����B��iG������cl���_{���^�7���6�Bj��u�O[?/98;?�� O�y�/����n/������ZV�*���~���7з$pا�6\��s�-����v��~��7��L��t��F~��t�yG������G[���:��>����x�������s�0.�%x�{V[�1������	���C�e���MПɃ�����w��n+=���m��v���R�y_8�/}pop������\]v��߲�<��ȟ�(|V|���/��r���	�����Z��Q2}������^����O���0��Y����������z��y�c��s��ǻ�^.��4[��k������7>wC}����	]��&�|�g��lD�\Ra;�:.�/�Q�>�>v>(�Y�[�|����qV[�eB�pY��l�}r�9Ι�7�w��ρ��`�b��y��?Y��5hwg��q����ŷ���e�V�cL?���I��|w���X�T��Wxt|��q�T��6����[�g����'�s�ߜ�/�/#���OW�)�|�.;�R>�E���!��O�C���ϲ����{�`��9�u���6ﻖ�	�Ҽ��N��O��������9~�-7�1.��n��[O������|�lީ��o������6��.���x�S+���l\fɉ�KQ/����L?s�"=��"���4��4n�R�6���m��e�S�������ҀՇ-y��_��-[�~}w2�͘����)�a�&R��%9 �I�E�k��؟��<O+�S������g��������|3�������=nC^��.p9���g�<k���,���k_�<��žWr�zY���0_��P>��|�sm�>������o��͗N���w�'�Ӳ���zn
�ש7f7����/�?Kzݝ6���
�u�[���ß�9v�i�A�uZ��I}����r>�Y遝���hC�0Ї�����U�bq��ƥy]pJP��O8@����.s�8�=g�����������ݑ�Y܃ǋ�_��ی���Nȕ��~��s?��G�:�J���[:UN<��}_w<��|�#���ܬ���A�Y��	%;�b�ָ:�?�i���⟳��6��Kv#��8�n�?s���y�x��6-oz���)��NxB�"8����Yд �����we��yo}^��?����%�����D���o����Oŏ�o���}�Y�S�	����|K��g��֟I;R>_�T<�硤��{oWmz?e9��%�����vַ.Wn3���g��Z&���»ǔ�(�s��sԻ�>ǣ��֟�����Lϰ����"���1�)��W�Wh��9&����q����.�sa}v9d���t_��=����f��E�����gb��C=����|�m�G�g�|����:��%<&����ֿ_��_Y�l��Z����uu���A���u������C��G�_����y�W��si��'���w�{����,ވ�eC���
_��8�\m$���EѸ\&��z��vr�7��Y�����t�bީ�8��ߴ�,y���*�\�����oT�~����p��<��7��f�r;��Q�k9n���|��;>��q���w@k���B�4)�x�ODr��o�l8��{�o�Oָ�]p�G�=H���-�'�O�o��P�G�bCo��:��o�{���$�o�����	�.��|w����Ӄ�u]�T��O�p_�<��1���wZ�e�]�����I>�5�	|���B�.
p�ѳ��;�����Ρ˾dW���}Qӏ+�rJk����mg��zKR�;��5�/���㾆�,>Ɇ�83�?d�����W2�å������s�</�N�Cn��O�s��n�uc��=W�Ӽ���1�g_'E������D�㘝�����?������i�®g��⨻l:N���1?A����Q��^T��&G�!��k���wj��lp�nm~�:�}��l=�66[,'��e�
K�xV=�h�8�O��/�o��@N�������i����"���W���{�y��?��3T>\R�:�ɡ�Q2;h�1�^dq�l繬��&��T?$�7�qG�r9��M:_��<����Wl=����G��uO���!����>�1z�û���T?�\�)έ�]'E�/��E�]�/��uֹ�::��U�q>Z��9�6MO�'�ZF������_���\�|����ی�־+��=*'��+�a�~�M�A�(ʟ����Î�����gz W�7҉�����"���c��)��4�����_��:(�c�0��/�����~6O39D>m���+`����ؼ���1�yݖ�y�'�_�k:�����Ԅ�7��ﳡ>�u��s9�s�f��vG���Op��sz�~��
��r�P�������h���7��#�������w~|9������s�ׄ������0���kt�I&�N������p��"��
��<o��R���R�h�O�Y�]$�Q�}+�O��ٺO�:}l����p����(o~O��ǅ�
���K���������n��3}��+q�m,߷��":�8CD?��3��������
~��?�[�.Py��1<[���p��Q��R�o}_*��}��}���<Ѧ�x����mxnE�)c�cپFϜeޒW��3:��yf��78?3��چ��n�|�tG��g�>�������/�ؾd�%���,����<�����k��=.�~���8��J�����Z���(��*=[8�!��������򪀞����lX��v,.��:���vy�tDq��%���g��2_�U������y����jw��g�1�.d�x��%=���z���^)��Uv�@�:���?��Gi��T?>�����q�%�W����3fx�,��C�5��8�.�4�M�d��]���C?+�½]��0�zu�����@�s�Z�+A7��?Y�mz��4�-���v�3m8�Y�
��9�������|�)�{gUZ�>���u���/-�8��ZL�(:����>��:Z�I��ч�y����vR�9_�ḳL(��3�q��6j�8��"��3�Y���0����3��P}�a���f��f~i+��|G�_7�Ǌ\uo*������
�<��:�Ů���8�=�\6"]�*�����z�s~P_��4*/�7rv�k������m��x]�?�>ߚ�1���l�-Qʘ�3g�{�?s>U��2���������!���K�'�_����.���_�%��aw|_��dm�yw��8�'8��u9d9�]\�Xo���:���v��QT?¿`mz5������������Yv�G��-U�S�'6�'�����p�ܳl�?[<O;�λ�����`^ ���c3�m���ݿ��?��B�j�����WD?��c�9��Q/�c4��G>Χ�7��Q>��nD�����}��9m��L�����G�CO"���x��r=�����{�W��y4+6��!���I�l�"y��=D��W�=lx/A��m�)S���X���y,��g��UV�ű�dz��;�?e=���W�!����Ή�?޿hD�����v����㕭���d��h���}�r�]�'�<N��و�h��e"t�g���>#�3�Z_�9�wf�R���'3?p����]�o�L��=��E[�!���Y�s�� �I}�+y,��ᣂ�����?[���*��2.��z�a���w�&�������{�2���J����|���������}���M��=r�C.w=��}s�������n���sks��?��]���T<�`���A����A\�qG~��kO}�H��w��ݯ�}nD�E�泹��Ʀ�g�Ǣ~�>|J��{d"��>#�ڝm�vqO��o��V:���$�VyP���h]:[���Y�������1�y������W���!���xsүL�(�G*o�s�o��w��nv���ދ+N�}��e�}������l����{�/���QT�e|?��ؿ�y����\2?����
�31��G����|6�OC�Z���%��}.�����B��Ժ.�|^��k�,���,�g��^�l|3?D����B�"��IvX�X�����U���y����ة���F2�_ϝ���y=�:�� .������p�G=ߝ6����S�s��?T�H���XZ��2?�qS�M�_�M���}1���
�?(g�h�����;��7�0���6;_����<�L����7�������b�p�g~���u�ߔ��>���8��Y��uk旪]�>�~�+�,�xl�A��8���kC>�����u(�]����O�v��z|���L�;�7�dv�����,��t^U�l�����}_/�_������g8�m�3:��&I�&�q�˼��9���;���|�����eV��[2�G�r�G�)��}��l��/�~���|��@OF��o��T��ݕ��k<��V����?3~��H�8�Y6�W��>`� �o8��?������fqN_C���=�{�����B�*��T��>��	����=�WH`z�_����׈ٺ@�ѻ
�w[�?��g=����h�_�a�~�����\?�w��K�zY������ӛ*�$�����G_KO�ٹB�=6�<o�{#�	�.���D/��N;��4w:2����A�T�D��]��ft}t4�y��|f{�}|�s�O�ع�Wt������?�b�k��N����w��\��K���[�{�Ժ�G���-���x���綠��=�����˦���R�����z� ���E��%_��k�����։w�Y�"������-��xZ�9Q��#�8�z,[�e�f~ �f#9����s=���}��;k}��%�3��w��»�Ud�u�����C�/t���\?�'15����/,���#<��HoDtf뾭	�&�Q2=��h�!�K�s�c�۱�|FR��W��p}u6�!�<��H�������;�7���\^v4E�D�|�t}Qm����ZY&�p�/�����
��e�����7��7�u����>2����%�pR�u������s�p�����>�%��o���Wc�L޲�O�[k��:�|�
~�����?���T�l�{�M���y����.d����|�ϭ�a�'��wb�q9l���7���ֲ�nY�E����S�N��ߋ�{���N��V�����_�/�o�u��Z��<���؜��mI�A��ש�E�����	�[;'�y��[�>�Gs��퓢��t��D�����^#�G]���=��3�zL?����h���~a��rrc�g�;	������$����?:���O}��q�wn��{�M˿���)�K�SiT���cl��>l}΄��k|�|��<�u��	�,���T�=/�a	���B9��8��q�JN���/Z���ϻ/n���??ަ��p�0~�-�S��{\���y'�~�ÿ���}K	<Zw<���ڠ��c�������'�chc?�7'��h�����;Η�6�>�E�T�~�g��=�O|n��y:�O�u_��w�ˬ�\D�L�gz����{����2���5���T]���l�g8���$0��H�櫭���ޠ~W�qZ}�>��b9d~�RaO����m��<:��O/��?Q�N����?����<`m�w�7F�_�c�l���y�C~3��?��*�Y������v�SA����	��\P_���s���rr��r~�}��ˤ��%�ޏz�M���#�%�P��U���^T���N~���+�w��a�O��&����z����g������Q���g=�� �Y������|V��pa��>T��&��������g��COi���Lr���_��}�<��C�O�k��|Q�ϊgz��3��c��p��޽^��vK}~G��{���T�=L��Z<�J9�s7��z��z��㈧��k.-�(�ς9�~i�W�ߒ>7�������}5���ۭ߼��oڴ���U��������Yq*�#nvbR_����l�&�Q2�ߍ�;�������8F�D�l�u���znx4����~�����L��q�3��_� �Y�3m���BP_�{���z�u��ǲ�(�'��Ǳ{�3�,����D����w�^W�y	�q���Ge�,���(��`G�mZΣ�=
�)�S;�Hp�����S����5�gf���c��`��!�t����E㺨�j�`�=��r��#���Z<.*�����l߼�.��g��혞�m/#8�`Y���YK����;����]\�������?JfGT�K?;�;��{Efݻя|0���x^����Lo�o?CߵڗYq�<��s~?��Q�����-p��|��m���b}L�g<h�՟���v���w�/(�7�����n���z^|��E𬾗��FqW�'�6,j77*o�;>O?L�������/�;�.�/��R���H�)�u���uq�ۭ��=3�7�uЃ��p�G'�$�ot�X�%�GU�-�'�uЂ�Eo��w�v�o�P}���U��Cޞ����c������{g�+��q�����*���������#;��|?�	�q���}Pc��ٸ�Z'�����u� �!��++����B��,(|o�G���<x���A��T?�C׵�~�'Dv�}����1o�����˲�$��v3?��
_�8�O���$�a����d�_��P�Y��ғ���o�q�uPw]�������\����<�X|�c����j���1�W�{��~��?�Ѓ1뎉����������������`���G��+X�}�xey�J��s��ǒ#z�.!��O���=o�
�����B�X�+GՓ�=�Y��f��p͓YL�`����5�ϒs���-��s��y4�"����E<�p�:�+��1��X�Gd�?[/gy��sv�Q��i/��fqu�#���������M��[z8��-�^�c���ᠾ��N�m��/�`��~�C����q�<s�g�'��~�����Z����ڛ>(~��o�����l_`����O����l����������g��?I���z��
��w���Ͼ��ݏ���_��S���;�=���l�� p���7���C���l�#ʓ��ު��І�W���A��˃�a.��ܘ�����se9�?�����0����ۆ�qrK��F�S���<4�V#�?��a�_?��5��x|,�f���Gp��ib��a������m*��]Yiq�����V{�G}i���!5;��� �������� �y~F��l(W��]O�x��O��zE��O^F��X���/J�W>O8
�͌�����{��/�f��>�����Y-�;�c�{�b��,�תgܧq?���"�#�|�|C���=��@���B�u7�~���� �KBgv�l���}������r�[�'��8�+`>`=��E��aex��NW�>���n��3mz���lކ�;���mڕ6�?�*'>N�gO�a<�� ��eL��J����1<����?��u�7�_�h����<����>/�`9��o�������&p_�9�������yCy�q��4��w�㴻��{o���G�1����7-烀W�u/�p=/�{�O��7��I����������Z�B���<���9�0��-#<h[���r^��g��|��5���f�����֏3����X��,~��A�~^b��E�����~�,�`lݭv
t�}�f�~�ِG�{����u�g���B^���?�z�u����G���|�gC=pb���8������}���2Kn[�Z�W�<U���%�����vVX|��}�1��{��G�q���7�T�^��C�sȭ�C\nֽ��.��2�ͻ��g�-��f������/��i�?/��]��$p��nG�s��s<~/��K~���ٚM�<>���1ڷuz����㸯�\�}O7tZ�Gᐧ{~�c(�O|����~ݖ����T��2t��T>t�ͯ�ܺ����9ˣ��G
�|6��d�a]��[fvܒ��	=:�<##��?�uQ�d�r9�߭=��T�s�����猴�W��ax?��j���#��3�od�����N�c>�\�]����w^��gU�`��� ���������i1k���dq����MK��q<�U|��F�/$x6'x��b�a�-�����/��b���6��u~��F������ҫ�>5��N���'޷>�>��:�3���ߜ��	N��}�VK��v�����n��~�փ(�~tD'�A?.�y��̋��+�1~��U ���@y���L���>��C���{ ?z?�����?�>��lyD��,����/���Wn4�'������j���l�?fm�༨������y�w\�g��3�sͻ�r�1�e6���T�'�]���!�g���m�w��LD��>{��>]��z��7��e<ٺc�pL~]B��zQ?3�[�p���D���m[[��E��C���:�ޞ�7�<��k��6|���"����D���S�Wv>:���L~f�f��=�'��G��wz��zv�|���u� �8�վ�~fPm�_+j����W����l�Q2}�����:�n�]�t����gI��u��G\U���G|��o�0��g�W�ǋ�%�`<e.wS�݆�:km�~>7�q�+��{}A���d�r<6�Y,��wm�~4���\�F�7��;����Sl@���o�����r_y��鱇�>����ޖ��e��=����A}�o��m��}���������3[_p��z6�'��y��}bJ?J�`��}�M��ֿ��p�3��W��r?��ֿ��<�Wv_P���$��s� ����_�^���	�����A[?�v��>�+�cd��j��p��8^�����m���+	��{9��q�ⴑ���8#{�r�RᏳ���Nx�����yݧ���~D�'�s��y>`C�eywL�΋����wI���#>�^i=/y^���Q����މl=��g���[�gx�ޟ�g_r<��GD�~ �������� �8�_̻Y���������uBP?�+��r����|W���=���_�y���O���az��d�#82ӷ=(��Y���x�%�y���֧����u�'^';�B'���t�Nl���G��,���K�WA+�����������w�����6���>R�i�H���=W�`�_���k�w���*���5?����|��B�3�~�b�q���yQ�J�o���:���kZ����f����~h��]��;�u���<�-�����si�}
�?�Ɇ%�/Y�.��t\n�����C�ҫ�nF'�)�S�*Y�~���Y.!�_�]����΍̋����d��]��}�����7*�Y���=������\��-�(�g�{x>_����/^d���f���}�~��}���_�	�7h��f�1F�����ϳ���sz�.�9�����.�������9_eV�[$��O���ak��	�+	�V�|��,��{{<�P�q��.��dz`�}d>d���KǓ�_&�����
�}=�?g��9��N��j�������g��R���휿���1��ׇ�N�(O���?{.�ۣU�W���m��u>K�L"�x���;>9o?��!�'C�u���W-��~G����y����+��\y����ԛ�>��g|��n�4��3;�{��|�^���ē�8@�nU�zN���پ ӓ�uQ�u��7�ó8�3*�b�C�g����򩔞�|�Y����w��d��C�y;��g���2=�/Y�a<�����s�z�7q����x)~�e���˹�^X �Y�N��~�|~���/�C��������ŗx��ి�I��S�y��]�=k�������p~/R���R�l$>�pΛ!x����[�k�?�i9��U�t�O���5&p�K�lm�E�qU�W���H��J�	�x�!��T������j�W1��~퇔����ޟ��X��ē�~�|�Z�Y��ཷx?����o\�?�O�O���>2��z�xz?@����@��E�l]��@��e�zM�Û�Ai�o����^ֿ*?���x �Y�"�$����Q?��H�����N[���r���G�aR��Է���S�\�^�|�"�������9����="���x2�����8�V�B��8�r�뚖80��Ć��Bp�}r�����OQ���u�r�ޠ>�IѸ[P_�.<6�������a�n�K�q�c��u����Xnu�nt_����t]�P?�����-��1�+��w-_��������{���4�����/�gz2}���y����A�L�~���k���y��=����1���7Nl(��G���,�/�y�%�_�셾q,?D��R���o���n�W�W\�A}ĭ4o��a�9�鱤�������M�ב�?(�Hn5�$��_���H���b���/ȉ�c����}}�q�,~����hV�1�B ��F�_�_~��Ц���>���w�n�b:�_g��IҮ�����R=��cui��,��J��q�1��t~y��ϧh��~�F�|����:4�c̲�Q<jV��9"�R�q���������1���v��,�9���~���������x���(>�eL�d���#}�nŦ���sY�a�~��l]���5���/����es���n&�����Іz�ϩ=��5�y����7��c���t�=�;�d�����Q��9��&ߧ4o�έd�w�����er�cx|�3� =�}M�W�.;-��j��$����ԕ�v��~��?�mx�#*n�c<s�G�>���~��ٕ��	�c�!�����B�i~p��'��7�e}>��������&h�]_a�}��8�17�.3��#�J�������3:���.�~����#<Fދ�����6r��U��7�'�����P�}�h�&�y���5�9_ڨ���%^�r���\/1���a\�������Ħ���y��:��v���L����M~������d�}�v���wY/�����������3�ϝ���Y�������_7<&��Kv��I����i�˓��}6�?<��}�1�#���u�fqo���F�L��h�mT1�Ӻ�����z>:�\<�GDqo�R~��x����S~f�@_������s�k�ݘ_�߫�ey�/�8n���yF^�f���6��5+�F��y��Z[���η�q����kV�ʟl^gy(:/2�+����g��>Y ��Wy�� .��e��֧Y?38�7��E���>��r��v�>�p������������u����e��s��1�^�W���K���W:�v�~b�����8o��ѯe���E�"�� ��_�����s�����`$o���g��;�K�]����	ϗ��2��{'��5���e��q|#�w1�������O*��6�g�x�����^g~�c���!��-��I��m�c*��*u����t&��x�vɦ�V��Kk�9Λ�8�aR��������Y��y��:��>Æ~��8Ugܑ�݇�o�a�uz+�7r���V���T(��k�>gy^��$��&�=��*��~�=E��������m\N�g�{2���ǹb:�qo.l�Ӏ����QZ����n_�_������7n�j���k�x�כ(��H-z2�/��Ggx�[@n[�,���կ%����X���9�o��� �����ǿYo����������D��'�	|�|��O6�&p�cD�񉴋�z�꫼��>{����Y�h����a<.��6]>;����y��y��?G��Z��|��)��w[o�^���J�l훯A��O
�o�۱���Q�d��Ɓ�?eC;���X�_��<��{����ЇHO2~���׿�����vz�U~&���~3�C��4�>����I���}T~��g=���!\��5Ѽ�}+�}{����~%q�9�����Ӻ�~u��Vؚ1����(������m������&��?~�	��CJ�,���e�D=���f�o�/Y�T����6��H�����e�A�l�Nl�����X�Gស�?���;�����}��2R���;��]�g��F���6����/�w�_�y��	�����zD��:,���lJ�>��x9�X߹��k:+��;�p�G�,�����z�
�9�,�'�]�d�h�oX��|>���P�A�O?���0��e��v���{��^��=��dyڑ>�v�WU/���*'�{��|����	G�_x�����G@�����v|�������$��v�
�(���|%�'K�|��^,$p���s�5��ϧs}��c���w�<�/Ѳ%�{l�u�H�̦��?�2�\��]f�:E�U1�,�x�����;�G�~�C�����������n�����nfџ�H�f��"=���b�c�G����PT�?����_���M�����5���s�j����]ټ���j؎���9������R:9�ɕ�C��q��wD�5�QԞ��:���U���i|O/�k]��~���w/��:^��.�����U�'�[��\y96�<�[�nڝ��-�Z&��#^����[6�����}��8���{�f��st�W�0Y������T�~�������r���߀��q��Bv�ssO+�������p�<U��N���r����˕����<���{
�}"���5u����w�f�2��o|?-�����A}�� o�ϛ`�d�8�l�?�k��˟\�����$�h���F�'q�����rnP߆������[?W<>�~�E��p�g����;�K�$��(��=����y������C߫��J��^�=��'6�/�K9������+��#�X�_i���6`xWĹA_�e�*��N.���=��F�r8�;#��l��m�C�e��X��k�������� �����z��Γ�xi�o+����h�ow���%�[vֶ]?��Q9�Va�
ܒ��s}�4�>I�dq�Y�-b�����Q �*�L��M^wņr�X�>���\:�ʷ,O�%T/�3���`��w�տ�w�v9{�X�G���e����akgeGۅ?���d�����_>'��v0k�ey���X���ݞ��Y�fI}K�GvpV�N����2���!��un�W<|ޡe_�㿠���Y�5��]�����v�R=�v����p=��Ɵ�.ӿj���������	�)\�_X/g��Z�1��V��(Φq��6z�q���R�C��i��z'�_��=�hO�2������w�q*���<��|���~����#
	�L�d��ߋ�| :^X����/>�����z���_�i���;g�ᐵ�<Ï��C+�ü��������̿�G�/׶���W�R�<6.c~��w�GW<l��=k�.��~=��]�D���^�^�|���~�K�g��W��#>��n��p�g������vNI�Gx�}����C� }��?��q]�7�Ϸ�-�.�ki������k	���P2?����2�O�3�:�����ן=��s����m{���;�V����>\_�؃Ó���8�|a8��;U|�}e��!A}��>ի��u�Dp���<�Y?��A�}����'�����N���.�_����␪Ox\��o�u���%������<x���Mu��<C�v[��Ժ~�~q{�շ�7�ű��ǧ��(z.���]��G~��g���֕�yv�p���{������+_�Y������z��(�T���Y���ڧ���I��Yqr�cݸ��{H��X?W��M�s�Y�Λ�6=.Q���y#>^�ou^�c�����lZ~�sO�W���|-��Y~�F�Y��^�C�����1������}-�l��y���>�7���Y�x���� =�Ær��K�OGb8�#��]gkq��ʿ���.ǈkDq�Yq��ϝ��.h>d&oY~�<c^�K�T=����/{OV�g2yh�'E�}�|����{dt�_��c���^��Sρri�O�۬<����d�ω�V�8�{y��g9a>�nq^�X��<KFq3]�^X�9<ҟ�ߟ�����{#��;g|S:aw!|8��c��g���v\Z�_+*��7�n�wvc��r�������.��Q���mW�d�Y������z����u��\Z�k�(���j���:�����|{߯������|���/��F�gZ��xy~����Z����h�+�����|槵��ϣ�βG����b������������A}իc�Z����x��_%�+�C�^�7fz@�~�>c���d�l�/��	���lq��(��\�����ϯ��#����������p:~�o�>U��f�Who��z�OF?Π3��_����1YN���I}^�F�Ƀ��[�l�?c���>��N�5N�Wm���v�iaz�����R����?Z��_O��z{�y���d����|�^f~��B|�h�q?�������Fr~>J�~�~����I�+��{�"�W�}�㾋I�G�#/�4��U��>&��
��A�v�,[~�j�? zp��\1��������o�^��%ί0��g�0�����t6�Q�_i�~�	�1�G�_��0����?�:+�''[O�Ľ��s�����/��O�ϾW��mB�|�_8���b����Ê������7�98�5���V�9D�s�Lf��v1�ϲ����R�q�O�T��K��"�~�֍�f~Bć(������ޯ��F� ����>�����ڋ�������ҟ�Z��[	�o4>���w��ܥ�'�/�/��ޤ9��|��N����p�n���@��;�s�k�7-������������?��>����������<�}����T�����9<^l/Xd���Z�<O�/e~��8�����B���ʏ���|��z���u\ ?�9�l�]�;�ϴƅ2;����9��D�K+�@Eџ���y�>Y+�#X�^t�xL~2<��D���e��O3y��dC~�?w���F��ˊ��;l���Gp̫��֬_?�Y��g���+�"��M����Q���~�ރ~��|l}o���8���9�����z����e�r������)��=xf벯p/��ݞ�]�[f�~9On��c9_��3�3\Y<*�o�u�Q/�������y����]�������x3?���,�����|[&x�~�s��>W;�����g���'���aWt���^�R���|�-hW�D��Z<�׼q��|����y�]��Կl��>���Q�����Q���4?O���N�r�'[�������s+��c�,ٰDtF������ٴ�\q~G~�Y<����1���p��N�)�[��Y�Ӭ]�����k��3�������e��D�R�k�~~y���T�����6/̻�8<���r=���]��������r���q:Ϸu������=�5�ߎ��~B�1������w�Y�_��[��k�_/���U���	]�Lj�˂v�?�'xԯV�������{�6�λc<e=��ݎ~���݃��[m�~ӎ�5�)G�G��s��o:�O�����2}�Mˏ��W�O~�|N-j���E������|�֏Y����ia�����~o����5v��m�{��?g���g@Q�d�>�|��ޞ�_�+�Q4>��ɒ�*g��[�/�/��u֯[%���v���{��K�!zne���%{O�����d8�Ǹ�����EdG����"���.�y��`;?G�;̇�uM������A�Ǒ�ش�l��D�g�W���w�eD�, kc�k�~� ���q��y��|�����Et~��@��{k=ǷBp�#�}��ِ���s�����o���/���Ag�kg|h�Wȯ8�6���v*;���l=�E���?�{f�%�����$�f�����z������#Ƹ�=zJ����Y���y�tGt�~(�����z�d�Y����=S�Y|>N��m�]��>�u����sGC}��p�%�}�Y�F�y|}-�gWm��-�����-��Dv�5E�s=���Hp�?f����3�3RG���2�1@C�?�+�Rm��� �]�����pc�G�|'��/�j�P>E��?>������(n0�`���ޗ��\9_�|,���;��J����}&�O�����R��}����Cޞ�Q�
�h~�λ�W^�<����y�"��=+~��?�����ue�g������{x@O�0�K�~��PЮʏ��O��*�}�V�?-xPt\ ��X�/�����]�n�6Z�����O��S�>�un�w�����G?[��c�+ſ���/�߲�8>�\��>�l�������WG��Q��w��/
������q������v�7�=�Y<���u~�љ�W9���a���'dy��k���H>��}w�M�G�9,����D|�h+������>�C��6�猟���gV���צ�����1�?���#��i����V�������f[�]Ey�x����K��=9O,�V~�F�p�u����-���y��:���b��EvV�|t��#���
s��uʊ��}����~��ϗ��)��X�N ��O$8��dz ;�	{�y�ȓ��ra?��wX�<J�����݁�_~o8���$������&��G�A��ϳ���O�kv��A}��Pf��F��.��.��oa'\Ƴx{�A7���������8��3��X�d�&�w(����Za��_Y����o��x)�'U��>M�j}����K�E��Ξ��Ǉ����7����={�zeV�������	y�{䥶ҩ��X�Wm�g��	�*�c�o7������WT����w����ǮûW6���-���$տ��u9��}J�?�u[��_��=�?X?���S�M�[ ���������@Lp��~�)�n'��iQ|��|���]�o��g��3��v�{����rA��C�Q~�^��K�O�:.�G,ݰ_^T�����|��=�.�{����&p~:�'>��W�'�&�aw�	�Z|���}+��v���>[�_cq�C���?Y��u]�r�R�ǋ������ߌ�_���~�E���A<�K��ظ`�d�8�'�w��a~Dx��[~nk�����1��f�\����=Xi��U3<��)�1�U_�����/Z��[
	�?3�!g��ؐ�������R�|��?��u�:zυ��|`x���^�{�3�\�v;�#}���襨��#;�X���1�7�o�
=�����LOg���������g::����9�&}�E��og����Oޫ�=�O���v��w�������Խ;�W'�|r�Gv����Ǽ�>���V=�D���u.~�ݯk��9X�W,�[�-���f�^��"z����u}���]��y�Y|#j7�gW:q^�u���]���u~]\�i����\?��'��[��S9���={DA�e���Y��#9���%p<�9)�M��Nο�~H�7�_�w�ǘ�ؿs��~ч��~E��8���=�-z%��A~���
~.��9�g�������~��_/��U��1�w;w=\�H���z���6���򲊟�6�߽`�p�]�+�ѽ�����^K������\��k��^�Ηl|u]|~��2�P2�i���}w������`�-�Sl�>�罴�+�]_�'�{�6/�5�"<����\,�sS�9[?f�\����ۖ��3<[�ܻ>/'�������#PZקT?ʫ��e����\��i>jF?�^3?'e����w�D�u�%�Ѽ��zg��G~�I}�ۉ֧������j4/f������W���w�O���9N��.˿��a��q�9�������y�+��q�;�����0Z���W�z��a��?-�iyؕУ�'[Gl��9�����y���D�z��-Q<x��%���&�/]�f},�q4>����8L�~����<�bC�-Ï��4�SY>���ɡ�������~���]v>(:��dC;��|T{�%�7���G���C�ּ_�@�!����0O.�W��qo�K�~�}����(�:�a>'��zZ��lײu���I2y�E�,n�g^�l���b�����6�OF�Q2�A��v�疿���~&Ϫ���p�>�p���Of�x�c\����'��Τ>m����?{��N��?��/���.Sgx�N�{���x�=�Cz�ٴ���>/�ϳp}�����!������w��2y�qa;5���?[D��ޡ�V�~W�����_�E�"=��֦W�̙� ��9�e^d���vM�S�gz{Ś�?O��Y�8�~�[N�|�+��I����8�>�����2�����q\�<����clv<��/\��Z~������Y}.ѹ�ȟ4���곏'����揯ݝ��?�Ær�C6}��=^HotQa~��F��|�����#������{�y��;eq����G��<*o�;�}����Skw�CQ9I�+���we�v�6=.�_���l(o���;l�Y�u5��b܌_�����߽����>[W�x��>�^���#��|!�[�[Q@�X��i���N��f���%z��E������7�/�'w�ښ�[L�G�g����W�g|ø��>�����;�o��ݮ����7tF�Φ��|d���;O��{��q�������?����p����R�/���Y�y��i[��7}�z}�0��_��\w~Ά��;�w'�[��2�L?֏'	<�/��;x]��
�H������&?39�\�_�3(�|�vqO��g>�	?��@�<�z��s?�_�_�m��~_��x������i�����(oG��w�}�|�VH�����b��+���>���"y��o�|������������� �ғ��콫(ٺC�U|���s?⊠�E�����p�dt��>t��[�3�K�ܺ����|���w{�l��������]ϛw���]4�̆��q0~�K�:=/�
����q��L~�~����O(�^P@����Wl�?(c���S�t�������8n���n9�?�i8>^���Ll�Oz[�R�Ԁ���\}L��Jc�w���*?[�w�W��Xι>���o�l���%n�qE��<�������Wt���w�S��-��KEM~�L~��q�����Y^.�{��z��|n����N����l����N�y����%�ά_��������m���3ω6m�|�ζi9���y#c��u��7��"^e�x��6Ю��Ü��}��~�kX�i��։���>o�'�oRx�$��}ì_��Z�/�z�5�K����g7�����q��s���I}���ȋ���^	�o-rh�ټ <��y�9��^�q��p�GvV�w��l�~��e�:���8��K�ᇞR���zo��B����gU�����	�D믽R?�3�{`����}(���}�<%�����E��%��仱��S�p������?�𤄞�����_��t��MA}�?Y�#�jܾ��A�ҩzmk�֨~�����{�Wm��}���)��C�����G�:<�{����݅s��w�ֻ��z&Zo:ݛm���>��H�Q������5_^qE��(��|����5ޛ�,Mc��`��܆����:��~2�';_��k�_���y}�s�Y�L�f��d��G|��!������/1~�۠q���xl}^���:��e�%O%�K���V�J��w���+�=�.o���&t���l���O�7�^��?���[��̚�x��^k��L��̍�gv.[�w�ڍ�!*=��#���ߧX�~1���(.m�<=���m��$����������)��{D�_?j�گ����� �����Q�+���(���}+.��W���)����������H�8��8C$������4��/gX��>O���my��X��^��D?�-|?Ofzܮ����|R@�D���Cez;��h����x��?����s��>���b�.��d�-/��E��}g����Q��S}�}w��申u��X�U�!nr��|Gα��懏�Gh\(�Cf�����\6�/m�^�������W�������g�g?��IW�k�&[�3e.���� ZG���h�l=�x���f��F�u۩�$���{�0��~�g���s���������g���3���@P_����3�R}�|�1���Y[�~F�q��jC}���+ף�O�č|��J���c�����|k^n�/ݫ��e�.k�K�?���=t5�+����o�v��a�~��:�~�~�+��/ E��'>?Ԇ���ڻ�}����N�+���wA���l^�dqo�8n��ϣ�J���:%Ó�Y�G��Q�R߻����_�y,��X����ߴ*�z/q~�O�3bc���*p����̷�+-��������W�}���dL���Ӕ?�����4ndD����bc~��4/���sO�����{ �����b��)���75�����A�7��E�×��Q5/�A������&�˿��si����j��T��g�Y�>���b=���<���Q~�[�nO_f�|���˫�-?����JØ_d���I}��f�g�ά�Yy#�H�]�w�\��!x�㼛����w�/�K�/�?�������[��yYG�lD���]g�O�m�>���r\���˘�y8o&6�O<\X����������J�{�A���q�q�8v�����Yc�m6U�;�>���i�{yt�9Φx�oy�+��F߫��	��#��(<{ϣ�G�����p;�2��[�饍��g��)?�<^m[���|�Ǭ��3�Ϙ�k�v|Q�l��d��-|��K�ȍr~��h��s�F�Uv�?�f�c�|.��^<��_��(WY�2�O���&p��d������\�<n�W��m��~_��W�/��@i�{������ˤ���T�	�������g�Q6Y�f<��Փ-�'(����]ϱ���3�/��9��~<+�ں�0������3	�h>?�!4n���~dtn���gV?[�:�1��x����d�����Z�^�� OfG���~�#��z陶nk��5ӳ������%��K�C�4Or�,��~^����e��R/��=ߺ��љ�#������C=/���m*�����޼��+�uf}V>#�1�Y��Ɲ�y�ޯ�?��E4�3�����:�ә�f����|�O�u�&k�o9�ٝ�,��:..GX�8��|ƽ(r�p�׈ʟW��n��{H�;��>�+<jg3y����M���s��5�t�_���o�߰}����\N��+�g�*��|���I�,�/�8\G��!\XO�����u�a�ߒ�Gϒ����+�$��s��D�w�4W��̜� ���� O��4����>��#Ǘ2���;��l�/��Z��m6-o�v+��b~���}�\�/H}�wE�-{_��Γ���s������l�v�q*���{�A��s��vy'�W�l8�9o*�g���6��η����_�nt�c�q<��M6�[>��tN��ў�'Y�a'���?��#�W������)~��ޣ�����y�!����ѱyTš�������%�/��Z��п�߷��Z�}��6-?�m��bg������s��x|�!�O�W����_��8b��=/��<����@��|?���s�3-��(�=�s��8��z��ˮ������뇖{]�<]�n������G���|���h�*[�l4��������[�=/��K6��x�s=KBϘ]sz�	����-6��7���#�$�Վd|�w/*��+Ku�3�R�G��Xޣ�o��Y<J����{���x^��k]/�>��Z��{�wx��G��a�_dG�&�'�?�7P������ܫ��?�W�yDܧ�]�o
zx��������w���������3�.�o-��Uֿ���3/�!��j�=b8d����l��s�$����v���E�ߧ��g��̟W��R�u��󪙟��#9i���b�t�˥�+�e�������ㅯ����2}��v�[<��uw��]F9/�1�+�M˕Ҥ�f�D��������{���EA�,�T���+m*�P��O蹅Ϙ�.ˬ�S��>��+��gz�7�o���g6N��?��F�7κ�4���֧�\<�.�η㤾����<�O���6�K�s�^�ÿ���z9C���f�Cζ|���ϛ��,_�%��M��e�M6�w1�SYiB�y]�|�Yi�Cp��z�`�߱x��k�^f�(�6�G��r#��O[���{\�(�����+��[�o���m��N����>�ذ�:��i~�������x��:�W*���>�{f��`��f�y��'�69����f�F��b�'��_���Q6/��k�m�	}��}F���;��N������=�'�6��8��<�����V�&�)�XNx_��*���[��#�s�Y~>���{z�v3�x�z�>_�����֧h+��9G0��q���������[�߿������|$���c���s���Q�V�"{o���^�;�]/�/���s��}_��s�W��f�<ld�������3��[��Vmxޭ�y�Cn3?�@����͆v��xe�������������|���6g>�������9�1a�8�����(�8fyh�zf��mۗ�§�����<�S����88N���
���o�ݍ�g�?��Sx�h̯F���n=�<V_�z�uD?�k����������;��h�&��@�+����c��՟�}��}=��Y���3[gEr������y��9KZ_��������kG�T9[i�����M˃�Ֆ�X�/ˣ�קi<�*���+��$��<��o"8�+�~��+]�����%_ȕ�3<}J�u6�7<g�řn���J�Y���~BR?�;�3��'��LFg�����(�R֎g<���x!��Q>��{��qB⹫�|����~G�����z���]��`2��*-��u�k��G�|f�w�����OFގ�N�(�����1�#ܗ�x.K�a<�s����U��8Ҫ���X!8�7�G���v��箞�P,�����=h���x��C�6�����C{z��Q�>��<��e6�7��Oc~�ѩ��疪����O%���߲~?�_	��S�x��>�}��{���}�yIλ�8m��`:��.�u!��߰.:_�-|��[���]�]���[�w��&��,�����3�9�ؚ>��:���/����������_�����d�Id׼�3�gq?�<�������G�y{r��F�Ğh4O�n����d����
����L�C�/xV?�C��
��+\�Y(���d�]�8���������M�!�ʏ�9��B�v����s��	�9P���� ��}ވ��=�g���r~�L����3��P�}����skզ�	~]���{�M�W��*��X���kS���>W��1Z�v���w��W�(��@�ƣ0O�����t�V-^���Ӂ=��;������s��I}ƃ��+p�o��=#��O�<@�+��'����$����y���+lz|�ϐ��~���ܧ�xn��g/�>{�M�'{��?�F�[��L?g�k�c�x��ǝ�Ū�����Ak�+�qw��U���r���}����y��c���~!����9�����r�/Ƚ��,����&\��^���}�s1\�Nc���y�Y}������,ٺ��𵵒���N�_�W���������f�7�=�|�Ot/4�P8�׌�ӓ���b�f9��j�3�U\�����m���I#~|��#�}����h�@��x}��h�Yvo��=�j���sA�����q/��V��6<?�tr����(ΐ��-6�{��L����y��|V?|�i�}ȑ_��q����r�����Np�'����
Ӽ;�����@�a~��{���Q����ۺNP�������:^x��Q���xȩ�%�[^8�E���#;��p��/��ó��,XN?�c�w�1{w4�h�i�#{4I�g~l��us������3���]�����u����Ѭ���~���Ӣ���=K�D�A�.�l����F|ݪ��<���ߕ��>�-=ٸ�v�ɏ�ȏ�yjI�l=��[��ο��~6�k?烱�sB�^�<"���:b��Wycy����nkvX��Z������;�)��������8����&�o���vq��4�����wK��y��l���G�{�3=�\a�?�����'֘>�"8�!}�Xvo���1��p�3��P�!����"_or�P?�\�p<|�
��#��l4�����+��ܜ߂�V������Y�4_�,�ҙ�C�2+?���|}Ƈ��ot�k|����-����>۩l^���S�Cȕ�se�:����B�Ãv[�E�x�|9R�w[۾�/�q��������X��LP?�2���2Ϸ�39�����Kk��Y,�^"�D�`��<�/�?��hS����
�y�Bp�"�l��_�e�m�%���]$�����9h��iV�������~ܢ��f�E�ny|��g��f��N��F�u*=�W�}O��F�Efg��Za���F ������{��=������p�o���1�{��,>����.�g��EqW��B�X��>���(:���'��'�g��~���+���3ǽ���w��ԇ��Xٿe��}�~���>���_���c�^�<��D�_�Kq��y�;��ҥ���9���L޸�<z���|nA�W�_e���}�+ꣴ�c����D�����l�I냎Lo+���g�m�&��Z����`�2��<��_�W��-�&����_��\�.��ٿ��;���g�OF�q	>���s2�����y?�E�t�h���!�'[G�1u�s6߳�	q��ާ�я��'��(Y<m��+���皏W>�\V�<��Ҧ���"o�M�%��d����.�����6�;�_W�	��G��ݝgCy;���~��F�eV���3<_�y�y��y�Y�ID��3�鷗�zg���r�y�}�}A��i�������]�x���>��¯��u�S���� ��u���;�k3:����E�TzN"���|�w��D������\���{ם�pߜ��~�5��q�Z���g�E�B�/�8��Wć,>�p>w�g�p�o�G˵c��o�O��u�f�H�{�Z�^v�Y���>D����ۍ�1�;���/�W^e��2�x\����c�r�?����2�! '�_�����D�JF��{�TnYol��/~F�}Y���yp�������?��-��п���>�~^�������y����,�������������7��
�y��szP�(����&��{�����6=�Y�Y�'	^h����ˬ��>%��s�گy۸�����u|W��.S�$�2~�_�g,y����N�O�����=������ak��Y�Ѥ���vWXv?��2���sl=���4�%�	�K˺E�_���{xTnU�g��?�z/�[̫�֦g��[	���<�ox=�1�*]Q\e�?D9�b�:����}�9���Uz�P��c�x�96�}D�#��4�~���~6.���\�uhf���(���v�]q�Ov��>�KXW)\�]�Տ���[8�G�w������r����J?��.5������H����	�ٵI�er��Q��/��{����J�Ё*�Y^S�n֯l�ܺ>�y���o�}���Dt2o �^�}y�g��{k�k-���֛�W��2�ڵ'W�ہG�[��}�ٹ �=,'�0����G(�����O���)x���i��0Z	���r�M����wc���ֿ��{�O��.-�	���H�����qc�ho��*�a�M�|���(�:���%�K`\��>�$��.����|8��F�1��[˟}e������:!���x~�j�?�g�8�5������,o�5^���~�8ߥ�����/<�j=�;�{�΅���"j�Z@E�l��[T�ў�o�/(Y���{	Z��7��̊s2|N~�v�}#����{�\?��~�|8��=�o�?��_�ǜW�����m$����Dv3�l^��B8"z̦�b`Y�3��N����{6��m2<�QZ������W��,'<�-xP�o��1�c(�ާő���W�}���ن�Pc���'��.��}nP_�['D'�m��g����{�l��xZ�9b��w|��pP_����k�#;��ex��%�?�>ifGά��X^-��M��x��z����>��C_=��M�w����!��:����l(�����q��}����
��x���;˯/�WY�^�l?K�Kwg����e,�}������0*��3�I4�~i�������B�yf�����?����_}� ~~��L�>DQ�A^��BgG�Y>�%x ��B�m�����[�S�)�[���xx���@?���'�/��M�����3��*'8���y�/��~���_����Z���+y�%�����𳝚O����a<�(���]��ܗ��^Jp�M~�|^��������?y��Zۻ͆�y��n��s�~Z������}��Y?�K�S*4��o�����l���~��lm���_��w�/|���G������}C��>o���Fk���=��s��z�>D���dtrlT���I�Yr��1���5����s"�����!���o��v��{�߯���e�%�g��������������f�rD஗wVz�:�~����q�u�U6<?���/�S���������jP?[w�8�7���-v���3޿S������iA}|���>8�.�������
�O�v�u1���-Z*?1��خ������|����fp�e=�~ՏZ/�lG&�]��\�懣6�FY�����)S��'ļ��I�o�3އ��tV���#�O��������Uw��;��?�����!'�X����y��|g��e�O�3x��[�]f/@������u��Ý�rQP���'�p�_c��2<�>����X�g��~������;��.�o�~1����>^gڴ�7�Ö2�w�vQ?���N������>�J��@i�/�go�'�vNP�S<gq����ғ�K�u�rb�z�:���+wVz���%�7t^�T�s���\F�W��3����'''t���Q6�/��(���|$����;�ؐ?���� �տO�~Mj}�7�';+\����u�1���n�
��>{�߿z^����x2�j�|���\i��&��]�?:�o ���G�������瑹>�#�}/����x8���}~��qTz��|������:�5~���N!x�����/pA_�)�Ug�1�)>lֿK_?1闶��P��<���	�I�qƏ���_�M�Ļ�h��Y��.3���=؆r��ʧJ��W�q���1����5�Y�}��7Ň�uAf7�<z?�?�H}�F��c�����/7��ߣ�'�n����W/\@�+�K,G�����A+�~�<~�|��F�ފv������]=��9O#x�ٝ�f�����گ�6��������g����Ip�s�wŷ�q�M���s��6K��\���|�i��ŏ��T�e�����k<z6E�Kg�=Q�:�V��16\/|����7�4��G�,�گ���s�:�2����x�����{u�q�e[���"���?�tgA��藞o�$�ra�zU�����d������?0�q?���-��)��u\�nd7Վg��}��uݥzE�I��n+׭��0.7�_<x��,��2.ݟ������ۧ�@��e�\j��;�5>�_p�C��)Mp8����~���7jg��gP��Iv��3�N�z�۸�s�����߬��M�G�O�tF�����z�5΃�2�s=��)���{���9�v��yv0��Q>ld�Q�U�g[�Y����~6����[�g��t��F�c���:����\"zZ���|\o�0-Q��'�<�{y!�Q��?S}�����O=���c���������ɠ�Y�M8�����[mM�v���3�-�In�%���B��q����A�/��Zm���\l��j�l_f�O��x��=����q�1=ܚ���G,��"�'w���~�����@?��Q:3<1��Pv_���M}�O����y������5�d�a���h�<՗|x_C�u��ҙ��5����D�p���	���x�~ܟ���7�X�ĺ������*h�n]���ڸ�oTN>U�=��_���-q��ݮ��7�E���7�)��UϠ���Ӹʤ��s廒���]�����G~�dyv>8���}臿q��������/���zv��\O�g�Z��q�M�K+�y~����K_�����W�7��	���
��U����pCևU���9���b8��?��ѾI�}G=��}������ۺ���ҟ�>��������w��寂�(���h}�w�Ex,��<���ד��ѣ�8&�G�s+c�f��tT'�_��E����}%��gpΧ�q��z{���ߓ����+,.k�n�v��;���ωp�,.:�Q~^c�N�{NP�u��~:�q�G߳���(~N�����kC=sI���(8o
t,Y��8�=��վg���>O����a��r��6-�vpL��Z_DzO�
�=.���q�0��#����>��y7O'�j�����/��=��2R�7�����^�����#�/�-(]o�~��ȯ@Q�N�';��U>ߑ�W��l:q+��d����h������,~��C�4���l�hqO���������st�\>�(����/4/��yL�ߢ�Q�;)߰�k������9�>�Fx̆r�v0:ǧ�hY|5��!Oz_\˺��	�k���Ӧ��G~~�� t���[	�U>�d�W(?}����������q��id{
����|`8�5�����?�>6�{������\�<�L2��=��)����E����)x��/������gk�oq��/��e�7��H��1,:�����?���g��_��z{q!��'�ܸ������$i7�'ۏ�����a<{�O�Riy�}}�-��I���Y<^&����aZ�lY|��gvp!�gq�l��J'���'��~�^�G����G��ϕ��k��������������G���,������|e���,���ϴp}~��[!.p���y�|h_o��az�\[DG����K_R�^i}�Q��+�&֯T>���#a�1��|i_[yN��c�{a�/�������j�Y���vg����P�8������E	=�r��������Ln7'��⇷�O7�W�K�J?������,����6̫�[�~�������e�}
��8� ~`7V	%[h�<g���z����u����Ϥ>/��a#zt��<��e�H�t�qa8�'\`���9k>2��%.�xV<Y�Z���&I}��;�;��_`����r�|��c�W�t.$p>g��d�z^p�`�{ĺ��m���_����znX�g���ze�t������j�������>=�~��{����Fn��߳�X�~+]A�d�Ԟv��#�}Γa:Qt��j}v;���������]�s���g!�m(�^����>��f�ޢ1?�U�gp�~����=���Z������g�o�����~�_<po�����,o\������C�}Ak:o���V�?�|�>e�s�����x<��(�O�ѷ�㬸�V��W�f������f���_æ1��q������A�X;Ez^�A?u|��4�_�'6<��c��}�_$�ێwX�q�!�5N���c;ŵT�r��Pޟ2�/e�6vO����=?������A��G���	�㕮+˸t���!:��6T��a���E��Y\��x�oJ�(��~,�[o�<d�S��vaO��/ȉڣ���9����̣�e���Y|o�>�$�M�~����3v~J�
%�����ۉ?�5}��Xn։n���!���^8�3]��^��l�}|���V���'Z?�7�l^h��_����w���e]7������鷬��Y��wՏ�`�z�u>������~���Q�X?�����g�<�M6��ȡ��?��=f���|fq�lA�ʭ��ik����/Ń���g�:��x ��{e5����Y|^^鹽>k�߮|�U�v_k�w�����װ��x&�^_#_A��D[߫>l��պ��������=q���v��a����5�ޯ��)���W;�Wq��9<ZW#�쾣���7_����h��u�.�뻜�.�q����6�6y�y �����叡h����oZ�����u$��dz�!��Q��|OB�G�����nm��s	����i�
��$���IR_�伯l^�>�����7����w������������U�y�^j��>�>R��+>��3�7�%������;�P,O��o��
�X@t/w�����c�K W4_�lZ�7Y�y%.,��G8>��Fp��z=^����%�'�#�w2����o�x��H<�������7X��s�8����j��b/<.ȇ�e�=WL�����~��Y~u˾6�o��d�����p��g~8��9�'����?�Uo�a���[KY~N���z��.m��/�;���l���,�َ��`���������t�������wGlz�<�l=���!3���M������w�x}�ӆ��z}��ؼ���������~N�c �3�Dp����x9�U�?�����?�xݶs�?��;�<.�� �ʹ��u��.�Ø/����covL�h��o���h�Z֗so#�X���/�;.W��>��U�c<�Y|.~�b9����}�l�P�8L6O[㥸�iنzo,R��}�g\ֶRţ����ݦ߷�������p��qg=��">�|���������S+�R����,���D������F|?�1����l|3?-[�x�~�}އ��,�忋��6��q,Φp���=�{o�8� G��Bg����?�o����[ʿ�y����/��e��c�����X�N�{�M�yn��Yk����<�=8b���ϭ#�1�~!��ۿ:����cm(��+��������qz��:���r���O2���&�窾�
�:/^_0p���S:�o�O���A�]�������G�n�>f�����|_zK���;���u��.��ezuS����|���k߉��Q�����x��=h���*�&����1�gy,���ei������n�1;�}������k��7ٸ<�r}���%N��9N��_ωƚ�I���'�3˳e:x��މ�Q����}�[p�Ҙ?���|]�w��������D�{M�����,���u�E-�E����P�����U�s��p;�f�ej���^�e��~~���i��ߔ?��s6�����x}�0�~�j���Wt>E�g�އ������[lz}��^Vl�?|���T>|{��b����x�����ʃ�^��9��gT���!A}�x��~4��]`8����ly߯�~N\Ѓ�A���+����'�����L时������X�������*bRdt��G���
vB���x���Z�C�_��x�2�s�{��v'�F��2>d����y�8g����S�3d�38쵞9�~����|����{���M�gzp�c��\Q�g���ߣ�U�mz��-�K��71�vU�Z��[�*ϴ�8�C]�����[�����6�E�mׯ��~��̷�����%x�>~�{C��^��'ߗa;�Z៳�<1�Ov���a����z\���}�7��(�"�Ӻ��+��*���Π>~3�yt��E���g<�yw�/�"�u���?�}X��g��G��'�P~�����Y����W��Dp=������y�������u?fk��s�A�Y�W������ܫ���<��6|�L��������=ڝ���*�ￊ޳	^���_>���c`,�c�!������~����#B'��u�f��"X�n<��������V�Yu�p���{��~����{�<^�[j�N����YL�3�2�O���OP�
���M���u��eU��޿�۴n����� ����k��g�%ˋ�wc|�x�<B���3<(:_��n��=��M���=W��/��{��/�wfB'dxL&��|����׽���� ��Ҋ�f��{��f=�{h<�S��7��ߋ�ڻ�uDo��g�{X��e�gv�������Mֶq������t��?�u7hZ���[���֏��?����
�ʆ��>��o��Y<���ϩ����~�vY�"�39Y�������{ ��/��l�b��:5��3�l��ep�������y���Fy��]vh�<�(M����YP?:���n���?�v�_�W:=������c�/룹���+���U6�1�ǽ����L�����vƷV��x�<�<���G�jц�u^��1�xZk�J}F|����u�w/�<3����-�d��{�[�j_��ݺ���&�v����'��}��ŢuG�_i~����R�e��oQ��?i��%���`?��J�	E�Z(������|��~��C|��l=o6=�6��jb}����Op��-|�/n����_�<��e���c��z����{_�c�hoI�����u�����'���ۍ�s�~���]a*����-��U\/�����(��m�> �3�5�Ćr�U�y��
��/�����UT��<�9Ӗ<�Lx}�2_��z����$��.[�����ғ���o�<���d��y�_��k-�ۙ_�u��Ж�;|�|��+[��ܼ��6����#ڗ��l���}��z���~��AQ��ܟl����r�S�o��ݿ&xZ�m�Vo���� ���о���
q����l���Z���N�#_׿����y�Ό���Ϩ��g.��m��2.hC�)l�X���;ޯ��ZߞX��z�p����������$k�'g<c���G!n���h^�q�֘�A��7�p��m�geّ��}����猲��<�����y�߮����}��_��������cq�,fA��@�����?������~��a?��H��'������a� �2�[�f�g�z��/�5��/�	��Ɖ��<ǆr��R�mڭ�OG:�D�5	����ܻ>X�g;���I��t�}8Ϧ�M����16��������[�#���Q����-y\�a���CV�*'�[��%�_f�u���8�CZ����غ������u���m����P��W��δ��~�x���W�Ɨ�~��ޝ�xg�����Ϗ8���K����gfv���g8n<	��x������GU�� �IB�	r��p�Qޣ�G��R���o������c'Mp~QK�Ԓ����h}�x<�������G~����J��t�����Y|/��_��8#��7�g����=�d|v���b����-���ժWѮ�2�gi�b;�|��'ˋ�������k��;@p>���q����w�H�k������{������6�����ι����Ї�H�5ˎ0����<������y�x���'<`���-��}D�����.�+���d��^Z�#��d����G�,��V�y�<^��U���o��|�E,_��|^��_�9٭z��/k2�}u��H~m#����4F��Z�2|���_�Ө~�b�̠��#���,�l]Ӳ���_��|��?�WM�������)���,_���r�:����٪o��,��%���,����~4�*ϼ��\����y�Y�����|���q���/B��_6�W��Ù]P�����<f�_ z��;mȇ�]�;��^�-�)C��}.*˲�v�.0|>�s�x��}}s�����*���w����<��L��%�bB�Z��7
�x�ę;�{~ ��ruQ����uk�G����:_p������f6���"��Y��=�n��z�.�R�)�g�C�*W��$���~V�j��lݭ|�)ߍ�g��Y�J����(~��Ko������x8���=xB��3zZ�xn(��a{m��^I�}����?X�7��f�gr�����[�{����z�자�Rv�t���-�+Nx�[��S����̺�1����x�ÿq�g��+;71+�Hrrֻj]�w�^�E���D�R������*��/k��?^~raA�~�,���E�k�e�g�G����O���q��{%x�����ͅ���s�6����	K���w�g���1�{Ц�G�}�g���xe�0<�7�~F����#{����9ο��y���bk}/z�ϕ��z�������;�|��o�������;�{ߨ|Fq���Xr��Ho���;2=��Q�g�3��<���Ҳ>��y���NOlx^#�,[���2��/�� k�6J6_��+스~�=<^���O"8�ǲx��J�'���:���n�����zGK}�g�y����}M˶����c�e/�����g��8>��G�}����ҽ���Y�d�5��̟��o���ج|��|�?����"o�����lx��� �����ok���g���~��q��;�_�p�'�|���;��,'�G�g�����]{q��y���7|����|]��I�'�3�>���TX�g?��W����"�V?�����|����+�.�s>���t�;���eC�����|�HǑ��?�o �z5�}��yb?c~�z6�P��~s�n|���mZ��.�"�Y�*=Lt���C��D����ڵLg��N�o��
��Q%�GQ|��1~���?�׃��Ϭ|��v�^�����\/�,�;Wn%x��>�N��i�fx�x��6�o���P>�a�r��i1|�D��0�Ͼ�ү�`����m�|�7:�KA����'jaWT�.S���Jgw��T��XO�\e�m�y����� ��J��X����W��d�^2�#��}�[���m�s��n�c~�<D�]��;}����J�+�|k�GѸJ��o,`��f�|V?�u�gl������s_��r���qa�_^��oO�i>�]��Y��|�å�S>���q�`�����E�l����ۋ;X�q
��ȇQ�wtG�q����C��(|Q�g|���:.�_����_x_�롋����l񼞥��������Oٚl���<b�p�e]ٹ�̆��]_��>;��Y�{{ٯ��l�olݯ<��ѡ���g�{���=�.�-���g}�|F܏�u:~�z=�������������}&���칯%\W�i����<��[��.~x�jlܯ�[�_n�_e־RdO[�{6�ikc3��%���O�b�=��o_[q�iC}��;�.h7�7��^W���6���s���u}��~4������ ������1<�s��ij�џ������/�o"?��ǵ6��U�{���w�6�ߏ�ި�l��ϸyL�8���e.#{���?����>�#p>���M���P��/��Q��B*~�Q��غ&���.��"���Q~����8]N�<�oA���_�0�����
Ƿ�}��6<G����~��)�z~�{���E��CY|/��Z�q��cDr8'�1���	h����-��s�?Ʌ�s��Ζ����o�O#8����e�E~Q�f���O��#��~ ��G�-�H�2;�|�5���N��>��v��j�?d|��E�ȀK�p�M˛�{9���u#{���\o���G�6�L'���=_�}#{+��I�m��Y���v$����ʘ��1�O[oO�|b����<]�5k���cyS�:�1�s ���s��#������Ř~�g}��Y��C�?�nt=��'�y���[��x�&8��=��
�$tr��u�3�_���[m�_�p�{`�o��r5�<g����T�c�8_Y��~�/�s���l}�r_MW<�c�i�Λ+~�����7���-��Y��}'�����<sO,�;��9O������L���?�C��^��;�R���,�o�w�q��{�wq���l#��42ܟ]�]���7[/��4�n�_�'��^ok�`�V�v�B'�w��g��f���Y�p�\'���X�A�Y� ���>�sZ��/,o[�19���u�^�n��?��[,�]�+�I}���yG|n}���s>���zs�jF'���3�������u�&�^���F������D���o��ia8�_.�-q�Km=7���d����<A��YK����O��#���//��[��]�}���K<hp�In���|��յ���<�l��9�t������
��#�m&'��U^/D�[���{[�[iq���W=��À{�v�P/��OH}�;��c|��o>��<N&oc�Y���F�lxf��X}v~<��|�}��S���a���?�P�x]���42>W+\���O�B82���sK���|��W���6f�v��^��'~�����Z�����39��$���#^�j���n���ߝ!�����?ۚ<��=9���X��ר>���5����-.��q���/	��y��e��%�~�u��6���y}�����<��R�;dkq��׳Y������X��xZ���aV���d�<��~��^��ލėԎ�~G�/i�7�ד�y����Y�z���q��{�N�0燞�D�
�H�[m�LC��l��l��F�n���2���8`��o����¼٦�Q�@g�j�Q�d�S�(M����x1��]i)�������߯�Pޠ�����7���a���@@��k`��mȷ�w�����s�g�8�o-�;C����v�^���������*�ᗸ�b�t�z�������=�OvI}�ϱsC
G���(�-��Kj��D��{����������dq$�/8ޗ�����I����u��2p�<]��Οsz@Әxc%��?Ap��e�צ|��+�-��< p>�z~b���q{,���߱8����5��Ǽ?��g=��O��a?{�6-ٺ/�;��1����|�i��8�(n�~����{W��j=?��	��}���a|���=�8��ez\N��\K��Xo�g�Y6�q�!��������Y	��⨘�j��O�'�G�k_����e�����q}�������(�g�ݸ��^���.[/��<o�q��8���&9F���c���ՠ__�}q�<�1�t���m8^e-ֹM�l�{M�7��1������r\����;��ûb#�N�����Ǩ��zN���y�_��0�Cb�;8/��ɪ����Z?�'��}�g���?�y��	�����ߦ�7�?i]Wz������#���_ѽ�Y�����6�3�9��=�tbq�W�Ř�������vH��e��m�{����L���ڽ%߲?��[��)6��O�p�#�������}I����<�3K�����{>��������K�k��ޖ'�}E�K��a�y�/�O8��=�׹�?/�i�<�6��3+����{�Կ�������<���>��{���8 ǵ2<�|�Ť_-����x�
wz�ȧ���w�iCy~��uYs��K�Z�#�:n,n�xN.?�\���]�}z���DtN�;�o�qշ��B?�����=�>O}�k^J�O��}�z����g���+&���!|�o�!+�S�>9�#��?�|l�5-��l=&ت���{h���6��������*ˣ���'��/C��������I}�����#����kA�����{�[��A�,��?���q�;���6�/q��������ǰ����~���1��@��=�.?�k�l/�'\��?G��E�1�]�N�dy�����}�,?�"�1 �z��3|�����p�	����{m�K4�~s�}��<�>����0O�Z�E��g3z��@�%{�����L�����yv�y�.��3v�>�OƇ�)���+zo��[e�"~��f��u��C~���������^�l�����n�Z����?��!�W�*���/����S��;+~�×ڴ\� t�R�g�o7��R?��øMv��r��p��������w��ϖ?٦�%��qE��> �w�yV�p���Z��E��q�]�7��[�%8X���Ys�)��j���"J|�wƟLn1���?����y�������������7:_��Y���^W�p�_�w���/m�~��(��n����������}z��c�]��l1?�����.�g�]������ؚ/0��R��P}��w����e�m8ц�]��v��p�#�-������I�����/k�����G�P:/���ȟT����>�����ml�W��ܱ~e�n�8�Xc�a����%��+�3�9���b�T�Ь�N��f��UϠ��a?t0����{�y��~@�we��P}�~��}��}����������������^�2�q��yG�������Ͻ�.��S}�&�Ϩ�v���6=�߮�PNN�p�/ǫ��G���R�������p{��r�/��^���ǡ_�A��T�#�K��Q��к~�|D�ۘ�Ao�&�?]�s���#�mn�NxfѶ������-p���O���[.|�^����tB�-U=��>�߅��<��띓�>���<��od�Yx̾��u����W8���P~ �����a�rܬ'9�L�#���7آ�}
h�~��+�c1��Χ�㹫d�Zk���Ć��|>%����1��,I�\���f�k�+|�����P�?ߺ���{��������m�����r��L�?�y|O�a[�S��^2:���ss(_�<���u|��)�՟�7F�Q��v����+?)���
�S����?׆v��~��3Hʇ(~���ǅ6*�k��WZ+��k�s^j�Qt>�dq`���`�,�:�aA}���%��;�Ͼ�a��\��}P��w��<g�	�����+�|_����oih����L�G�w'�}�_���vu��8�?���}�J���u��1o�N�_�+�{f�g_���_�~}�r�����k-�X�/&pЯ~&��m�?�����z<�M�_�74� ���,=��l(���߆�����i�A����8��)���y����3�O�;^�[m�y��*����<�)�s,��q����=��s�<���T\��v3;����n��y�M����ً��h;�Gqo��B���}Zy���|�zH����
�_�a\�������q$꛵�[�9���˰���e�X�e�|6��~���5��bm��8k��o��n�~�Y;�2z��l]3���>����cW��^b��п0�c5og�}d{�:���I�x<��y��W9/�t�C����³s�<.�*���C����Z��1�c��<�����}L}����c>D�Ϣ�z2�k�|�ω�_8�rEG\wN������ѓ�O��t޹����g�]O�9�h^���������'���qJ��@��7U��>����lZ�T?,غ,�<B�J�Fx,�G�֨_(j����b���zO��m�/r�A�|�e�q�Ι�Ϯ'8��k�=]�y�:v�S��~�!��> �x����fm��/��۫6\G@F6��V����d��+�,�����x�?w�����g��b�����p}��J���q3�.��z��?��O��?Q璜����/��^e�q	ز1����,������=�W]����c�W�k�{�7�gj��u�dC~��z*��|�����l�����b�qԹٯ��Gcx��i��9��q'�����G���?���)�GT��lQ^�$�s���'�؈���]]>��^���������<��b_w-V��3��?���(�y����z�7������7���N|��:����� �y��e�l�xߐ���qu��X�k����pW��/�a?Pг��B�~��v����p���+x���:�!�O;[��W��2ܓ�9�=��g���#J�v������:�hb�y?��n��S��,��p��~�����M.۷տ��Ϳ��6֡�����ǭC��PT����+�7�N�ϭ��݇�su�_���zT�Kr}���*]��������޿���7��5��k'���6���`}�������0����w�_���s�·�x��v�z���n[�#u�_�P{����8����]Q�G|��?^ag�u^���-��%�ۨ<gp^oFp��,p���_����K���Cz����r�q��V}{e��M:S�m/Ц�T�ј?��K����v���Cf�52<F�#�:+*ڷ���j�������⸨�'�Z���+�MW�h�G�<d�����젾��ڧ�����B$�[l8.�<B��\���O�9?0�W�#��������!��	��A�N����ˡ�7�o�0���I�l�/�/�����вE���m*|�U�ss��<��:|�l��y�m����n�����_�l�I�Jf�2>h���{
<��7��|,}���A��~FO��fU�����п����<�v[��!�g�t|<���\u�O<���6�g�d��Sd�c������p���\��4e�<�ݵ�l��"q���3��(��ӆ�;����c������9N�2����}���@�� �� /�g��=����AOj��\�����>��a�#I��A��0���}�w��³�0�l�/�������|m�y�_W���	�l�k����ڦ����x{?�������U�������]�(�C��k�����qk|xw%p�?�XՓ��g��宒��U��qv��F�R�~�gPZ�g�����q<��R��}����/��k��_�x�Gc��q�h����#�P��_&x��������zX�gh��_�o�{G��u�΀�o�����u��^�kj=_����8s~&��-�� k>���{��6�w";G��������oX��q��^;/-�[���oG,γE�AϿ���
��/��������Ԇ���M����h?.���毮G�v���iد�LF�M�;^�a�
��O��s�;P�>Wv|9A� �v��GU�i�p�ӷZ��(����g�R���9^�����r������Qt^��0��
�31o
�X�#��]�7�>/�x0�8p�ʧ�v]�;�ϱ��^D&W��[�����v��3�Q���(��M�+}܆��X�k�����w"p�����&p.Y|��g�)0�0w"��������lD�K���E�נdz���Cy}�9+���[��Gw��5R�1��Će�7Ĺ�+�k=�?��c����}~]У|�}��<b=���>���B��uFp��Ǜ-�/�����Y�~�{���������Gc�ǹ�GJ��lY��v�����#���x��Wmz���=6��k����~�����8��{?�_R>e��>[;c��;ʟ�Gv�ƹ�s������R�J���q�uL�|λܗ1�����껜�,��V�߿�����
w��F��W>n��8�r�き��v�C��GO�n�-���'�r�'�I}͇w��\�'x�H��Z7�}����3��}~G���w�:��
���q9�;�,]s��BΫ	���f��x]������z���[	�U�������͋(�c8ǻ"�S�`իk�l|�нl=NE爻2N���0�cC�|O�sN�6?��Ы��>�ʹ�ګ�_wd�F���r���q��l<�r����9��<%���W�˃�?�������G�[?���X���=�|�Mp�_1�mXTg�S�s�e��F��f~�1��Qtߟ�Gp��e�q�?�����M�+��������W*���>��[]����3{{�y��Z��vgC��d�υ���v�u_ �}���}�����ؐ�����͓�v[��������
w���ek��P�� ���H���}jg�~�;�w�[���g�dz�~��u=�8�k��~����}`�vqA����7�OF����-�cW�����C~T�2=���=�ot����>�Ć~���w!�+�����w����5a����|��7;�w������w6�~��Lo��!
௬u=?��g�����L�8�|���ؾ��gS���>@�$��}OཏЉ��JB��ׇ��|f�c����غo�o�q��>d���_P���'����C6.\"������W�tFz��.�7Y�:h�&�ا[:QO㥾6����;nW�d�F�י�����&�W�w��\ xЮ�w��cvS�������|/.�/I}���ϗ,���t�9�,_�@�,��[����|?���f��}������;N��o��q�k���jl~)�,���Z?��p�q��ǅ ���x\_Nl��<U:/+_����T��y@^G�����N����;��ϗ?�m���>I�j=��S<������-���5����|JR�i�T�x_�m��x��^�s�1�+v�6]?��_.,�8O�v��ㆱWz2<��:�G'�3���;ǁ�]��6�H=�?c0�>V<�.�0�c��_p��/�㷀�Z�9=��4����jmzrldֺ��W�n�mM��Ӷ��{:POw|�������[6��/��'?��}T�ߺ��F�����S<c�̮���p��&A}�w����RaYޝ��^���?v�Y�>U���iP_�;���_��p�����6������hq\��{d�D���Ou~���<�	�/�w�^��m8^�ϗY>��Ǟ}������������'�����Z,�ټ��^xv��γ!�{����Aۭ�p�^�~��>U�����	��|���qH��Np�����l�?�'�E��-��� �N�+x��s��T��Z�=�W�=��|d�m]��~��pD�\��`�eyq^x�g��A�5���w��������{
c~��ۅ�������o}������|��Ax��j_����]+~>�Տ�;� ��ש�p���
�LU�؎d���Gf���< _����|o�	��?��3��zA���o8�o��?��l.[�T�fQԏ-u:��������>��x�V��p�ǯ�G�R��1�d?���~��6�����ڙހ�Ř4��~�z������a>���y��6�Q6-��M�Y��/������(�̱y��a�yL�����V?��[~?ș�O��t���J����g���q����v��J��Ϗ��	�7��_��uƇ}�9���X���wцr�<݉M��f��<�d�<G��~eq�̎XR������8���5��xc��d�	\�g~�����9/���n������wlz�N�x]���>��K�m���dC��{�������_A}��}Ǿ��S2<x/���f=��1�>>�=H���(�|�����e�S<�;R���}��m����df������g�Q��>&�ώqW{{p��3,���~#�/���~̡h����.W?d�m|D��lm��/�F���Yx@���q�->��D�A�黟�v������y��]�׺�\��]��Y��Oj}�.��'��̚�����#<���ƫ�>��|^���qd�:�α8ak\7���~�gx������ό�x�6��z8�[�N���4F�����A}���"���sf�e�S��`g�X,WZ�wW���q\��\q�.��lZ�f��<b��{x.��V|��"g�e���߿��6�;ۋ,��+1�R�Ӫ�9Z?�������>�����u���Gx�����6ԫ��܆v��
�)xV��{��@����~�|�g�<�|����'j�G�F�������p܈�sR�l�O��Wm�/���}������3�7�;�.��l�8����)�r�S�_�>;��g�Q\*W��]wUz2=?F�����s����������=چr��o��s~�m0^�L>[��\G�8�mE���Q<_�t�V��/�#>�x	�ys�'�o�]�_�(p�7[�7Z�_XG?T迦փ��xN��;�ֺ[��M���fy�Y܆�H�9��y��y�����1�C���+c8bQ�#��;mgW��98�/���M�d�n�4�=���L���w��P޲<�,cko��c+��P�C���K׏���}#��B�凸_�j���*o�����'�W*��<����;œ�O�`1ߴ_�(�|���6�?6�I���"�!��^V�p����zL����Z���;@p��������W�E�yv%����zaw��96�{9C�p|����;�#����,�A������8����srG�g�]]_{}�=��_l�.��?���F����y�,��]�u��|�d��w�c�oņ�9���v�}C��!��8ʆ�QԞ�.k>���X��]¬���C	�K	<�o�����9[��,�G�?�����������(�+��;�����X\�������CPT?��]���D�s�3�{ϲ����Ŧ����Z�?F�����l8�k�w��A�.�mՆ���������(�~"�Z��%m;�3�Ϥ�U������*�L��pY�{�2<��v��n$�<����">+�"��:X�߆��?�w���^��\��8��k����ջ��+�%x���={��(.L�N�����>O�������v}�!�5�C���z���_�~-���Ր�V����Wަ�e:ϸ������/)�~k�g!����>����y4l7y?�����}�[�ʇ���i�o��.Ɓ��c�^�� ���e.-��hi既d��̎����^t�O���ع��>ho���|�X?f�n����D��(\��9m�3��1�X�x�;/�w�~�9P��܍ҟՇu_���b�������SY����2�}��*��sR�����{�[w��cC~��W�z/��|����@t=5�:�c�߭������9��nOW����O����Ƕ��-��[q���~ue,v=��/�����xo���{��_[>l_|yl��.��:&ofm�.�#�#�������(p�V�þI�}�;�������}g�z���zr#t�=��7���+�ϳ>�yzk��1=����į���%���<��m����O�G��+����`]��b�p9�3�3*�,�1ۏh�ݏ8R���K��K���!Zgi|���2:���e�ӳyw���|��tvOZf��Jk| E��<�{v�.��\}��w𾤷�c���d���x�Ƭ�-�,ޕ���Ѹ4���Z\��U��k�������r?�H6_&R���#�O��y����X������O���?_���T�T��^�]/r��@Β~e�F#8ӿ9��z��L���<zϚ֟T�v��gk^��w#�b����]�}��Ĩ�|�ec��}c>/��j��_��*sl�K;�E�_��4k�[�p����ө��ǣ^a�;E�^D�]gT|��a?�� �~2��̯@�%ꁲ�]{Wơ��S���3���LN������O�}
g��e=��t}������E���ї1�����s��_L�0��_����)�=�b��r��Z����ݫRvm�5铮ؾ�O�׷�����'�Wo������y����2�:�O�4���Ѷ�'h�����6Է�������o�*W<�<�<,�q���#�8��P���J�����{��<�� ���<�c�qA<d���ZG���=��`8��19���>a�\l�������=,���o��(��i��v�Q����x|.�X��.t�ޯ����Mө���\]���	��p�s��_P��.�B�x6��z߉]�n��l�_��w���t�y'�3��H����<�<�P|�����ؓ�ߓ�����Z�E���#��{�mk�5x�#�Wg��	�.\Q�.'ѽ��
ؿ��7�����g�
�'پ0�/���{�{A�
�ߨ����
w9��_+=\��
�=��a�������	���cG�߿�{��5��+x���}��N��x>Y�o�8����q����x��wx���oX��V�u�%���w��Nއ�v;��G����_������zyyB������Q��o�,O����-�����k9'/)=��,/�����:�ʠ_�gܟ���ֽ/�S������@p��ϱ�����{z�Ï�t��ʧ4�%�C�qU���!�g�򠢸e�nw�����ϧx�q������s~/�6�D��s��4�/�S�Nlx/���ޯ|���_���_4���e8��g�'���x)��S;5k��dE��]E��ݧ�'��o�]��Y�?��=��.͇��E���qi���<���5�y�O/	��v0�3���i��=f�8�3�_��}���֟o��}�7�~��(�.旞����v��8?���s������v�|c���Ć�eA7���2[�=G�k�)��^�m��� �u1�7�͚σu���Gx2}�t��8"��u̞��&�tn��<����vuo����2���m����Gp�]X��
�k\�[?�~�����>��5��Q��o.�(ά�m����ζ-�lܙ~^_�~:�+�����>�g�r���Y�	w��z�ǌ�ù;�g�J������Q�]V	~}�����C�.�U�l���-��'��+���߯��!���f�W�T�g~r̯֯[�ϳ�b=��gv��}a��Y��O���������]��28~�ݪ0����w�L�����y�y����^���V�K�'��L:��;���?c}�ȿ��!d���߻�1���[�����v9jџ_�>����쎶{V}^-�#6.ό'�S��?��+>XPټ/�)�E���A�0�����=_����A�7��a4O	�nw�>�)p���<w�S��\*>`���o��󅠾�[��ϮG��;l�z���<�QTh|���`��v*���u݁}���(>��~��A���5��&��JO�'�'�f�j���_�F�V�9�k�"���v5>S��]��Z.�O�3����~�3*���7輂o��8��w��A}�1��D��wk�0�o�g,^4oq��F��_b?���L�y~��Y�������]���N���o8��q����u����;��������X��'T���#�xiɃ����9z?ʘ|��;l�o��g�7�#@�Gv��n���j��p�_�-3> �����~�5��Tx]�v��
����A�߃	������ƿ@����j�?��}�J&(�O�g����W�>�⇜�����y���&v������*?�})���5��T�qy�n�>]+�x����G�S�E�NJ���B'���G�:����<��;=�?���i����)=���vU�Ŀ�k��%��9|U}~���=r��yPQ~欸w���5�/��y�������=Vަ�ct�*���j�(�=���������}�����eXğ��3*��q�k��yqg:]g^f}���?�[K�<�-���s���z����;��������Ap��f���^��|!�)���~���{aԏ����s���w���{�w�ay�u"߯���"<4���ZL�٥���:����)�����~������A}����r�_��a=_��ڦ���<�?]���ͳ^zwm�,���N����۟���.v}�d�����W��}P�����×l=��������|-�/�.�����*�'�Ǽ�>���W<N�'V=���a[�}i�3�/�ن�(2.��5���<��fO ����s�_Z��&<�X�=��/��X�X�/��Ŏg��x�m�gz�{�P����	����y������f�C���'�^�
������G���W��eѽ^�گ��f����[�����+-��;�G���Dq�{Z���A�r�v��(N��������>���~�w��o�ܜ߹򻶶������#>k�uP����E��lG��������7�|��<ϸ�s�Y�������O�?�����[+؟9��i6���D���{���㻿��}ܳ�66�O5�7����O�5n����׬���o�����u_D����2��*�?�so��Tٍ�i4��m��O��|����<��C�/�d瑕��G���z��j����`��a��*z��?ͦǽ����������W;�q����#�c�엮Z�r����W+�2����@��޿�t�_=�����̯��k��~ߕ��Zqs��گ��-�\��L�A?��;�������Ug��'?W�~�|>M���������ݯ���ζ����������3N#����z��
��O�Q;��� ��U���a_}~��1_&6�/.����wd_�݋j����=)�)҇Y܌�����j}�a����M�Y�ž�������O���v�Ϛm�����ߧ1��u������s�z��z캠����}j�k��=��p��:���׆��6��"�������Yx.��ˍ�G ��� ��va��f�~�v��.U�O�k���g�
eA�|�����͋V:ѯLok��oz0���о`\O��?G�y�~^������� �p�������sY����ǋ}�F�������Tz�}��1P6����v����1H�oY�#��~��?�~����y�o?�_��o:���}�߱�����oc�a��κ��ߩ�C��Ć�%[�:��p<�}A|�;��Ӥ>��<(�3�'�+='R�~�	���R~B��t~���~���|6��?���� ��Y?vg�߽���9���<�~��ϳ���<�W~���8^]����͕���w�=�<{|��������~���s�m��y���=���w ����g�.�AQ��Q�]�2������z�M�W&oټP9|u}�}�'�M�gx�G.��_�[v�������z�W���~���x��/�����˙���_t�'����G5��e������і��z�s����>���Z��J�WϬp�1�'WT�����Tyf8�w�1�{�d�t!������-��?�|h��x���Ⱦ����]����A����a��ax���������}t��@6��	Y�?�~�M�)�)�]��l(�Y����������I}�og�����V}����9�F�E��:��=<��c����T����1~r�Xn=>��V��?���ZoN�C�j>�ؼ����ȾR�Wc����M��_i����Gו�6��-V���n2=��Ku�����h^t�p�e�n�����"آ�P,����_��A�ǀ?�j�����'�������4n>d�Y�����K�C� �a�'�߿��}�M{߯��.�ɕ��@����q��+������Ito���x�~�| _������u_��E��}^_��Y
ן/���z�6|�z�d}���j�x���Z�L����d�]��������Ft�m��)�����΋[j��߸?�q�������	���ek����c��q�_����߽����}Y(�\��#���c�W����תG��k�3����n9ϵ�>/�>D���Y����>&����"=����7��ﳟ�pK�~v��e}�tAP?��,���t���U�Y��Q�f���?�όŝ2�}�y8�����S��w�������~F��Cg0=ٽ^\XΗ+L߻���g|v��x�I}�K{���/
���p�ך�g�낞�^��+_*C{��E?��q�LΡ'UN�M���d���C�'X,?:�v$p�&�o+���1�f�M��ޣ˔�ݳ��ʇ�
;/��v�rdO@g�O2�~�|76�28��8�s��3��`z�?n���1���Q�:^��_�u���E����	~��:�>�8�M=4�	<�to���>vo���6��r�g��w�bO=�i�'lz|A��7��QA�l�N�\����O@k���6�w�}��ӝk��Ǿ}+?[�Uy�q����g��mN��\�sؿ��Ac�o��D�m�߹�o��Y�6۵�<�ˡ�F���s�= <��^���<{o':��tf��Ɗ��ߓ�y��5����?X����\��]֯��y�|��u}9Y�o���ՇJ��x��� ϼ�q�V���.'��\������0��x���w	�]�����^x��x��O�k�;+-�׶��p�*����,T��x���%�k�|3�W��*���c�6���~?�笗�"8���|�w_B��W�W}��,ާ��$��c�_��v$�o�:��?��d�̺;����8]���~�M˃�ő2}��:d��M����a�/�Y/��Ϲp?6z��P}غ���-��T����VD�+ߐW�x�����9��=��·�u��L��0Ζљ�9��g��벇X���x�����(���(��<�W�y��u�'�bB��æ㱼����w*��6}^�cv�O����8����m��=���1���
s}��_J�Jd#�5+nO~ݜ�}�y��U�~����y�z��6[�3=���p�g�4&�K�����F���J���[���Yv'�[��6[��6��}݇W���>���{#Q�n.W�iRx�Zn�ԟw���Y��Za�G9=����?�v��'mxʒ�wX?�^�!��塕ַ��b<|/֤��e����Y��R�Kd��4��R�t���i�vX�_�d�<��mQ�/��(�Z���lZ�b�ܒ���������8BN�N���u����������N��<��p]f�*���1���[��;�N	�+���S�u�[����8��r{�z��1���@���+�f�����5���fC9�u�c���{5[�5(j�ήkH��0��_�o��~4��<J�^6.��o�/��P�o�/��h�8.�X�c��e���G�/z�*��Y<��]a}����m8�������o�����;�o��&c�l�������\�w���ۆ~�1�g1hW��U֟���'p=��r�W��z���<�S<���m�ϱ�x�M�/��/���x����@����q^�����'��|���,=�p��}_sP_��¿�ڻ���T���	I��V��p?�3m���Ex���I��.�^���#�=g��6�xP����뵮w^��u.�t��1ÿj�,\iCy�������k�ys�/�4�w�̇�E���s�2�w_q���u۵*��b�P��\YWl��R�F��{a>���ι� �>�>�z���!�ݱv�O����s{�.���*~��=����A+=�e�m���yp�&�{پ[����H�!�S��^}�GE�����{^�D�T�%�K�7��_���n�x?�����_��~f&'�g����=W��>�+�}�Z�}+��^x������l�ν��s?��b��_�W�\>��u�U��}�������*�es�k	Z�3�g�_��u�Mˡ����}2��Ep�G�&��!o�wslq������>���;؏�{2[�5zfxf��u�ǩ�>��2���=�GY~O;���Tz�mA}�����ɕ���@���l�g�g��/�Ec��x���<���T�ϣ�8ߍaA���jOY�q}��Ϧ�(��G"���w����B���,�����ڻ3�>�ߎ�u�/���w���䑄?�L�#�����g2;⾤ϱ�����q]P�b�q{�ߦ�1�笼��3�Gr�Ն�s
�E~o�_�t��~w��r�Y�u]����N�����������I���I�؟���z��~pys�F��YޅY�h�K�y7��/?\��|�D��� ���O�c��G	=������n����M���+�̡�}S<��h�虵����~6߁G�!ے��1�_�g��|e!mg�c�V���g���t]��Cv^�%.=F���uV�'6�'[�f�dvP��I��a������<T��o�������Q;���z��x2=��[����.~�+��~���0��~|����	�]bn1&��������~!����,7�_�t��>he}������G�f�]�@�����|~�T-��.�3����=��u��Ο"8�`G���;�u�GYM����~���=A}�gܿ���/ �{�"��E�W\�O��7�wO����ӏ�ڙ�H�*~ǁ{ט�M#����|�8�/[��b�w�O�������"�e���W��w��Y�v��z�����i��ƅ�ޙ�4�����z��ӱ~��=Xn=n�1�U����xϪ�e�,���h��N��j}5���3�q]�������^d�E�᢭�y��3�G^��!Г�W��}���&6�ծ����+p��<�x���}(�(�	^�����W�t�z#�W�㜘�EW��|����Bj�X�x��ܜ��=�|���9��}F'�/�������_��0�n׾f��	��G����qA�T�Rx&?(��%�_�ֹj��]��0��Y~�#���{����U���,^�z�̒�.��9g��ã{A�>�z<Ó�y�b���gЇ1y@����w��q��ˇ���s�Q}�W����>l�xxHϼﳸ�[l|���^��6}N���"� ����<�"<��?VXYlf�����c=u|�G�ף;�I�2����\���M�Y����f4�wѡ������!"�bLo�^p�q���[�`��K�g�g�g���K���q��Ļ�������7a8���>��E���ˋ������V���w��u0���gӾ�����l�����(��G���V��|@���q[�1�ϫf��7������ܟ����3�U���3����}2�����	#>d�Yq��~���.�������Q=������86Ǉ����O���
�3���gml|��LW�=�>�8����%����뗳l(珨p�C�1�?1��?�r�������o�uOtom�>�A��~��+�K�>����f���M뙌~�I�,���3j��,����>.m�w�ߓ�}Η��7��~b��.���|�fx�u���d���XD�?��^��%�Z'���O����Y�O6�3�A��o�b��X������G��vƟ��{(�F�t@���/h܏��r�����ѽ��u�"�0�j��X�w���%v����|Hm��x/���������z�}Z��r.��|�/���'�(�Uh��'�ن�
�+����,�#q����y:�G��?U��\L{����׼/�OI��M����`�2ߺ�3���-���8�%�ۋR3�g���#�R��&�.'�U�h��Ctϧ���*џl����;���Vr���Y���N�;uo+�[�z^�!��V��p��������|~�D�@�ϳ�m��9�Q9��>��P�:�_�>?��j���o�.��l��N�3�y�����?��f;����`]�p�_B��������|^&��곏'�3��*�����Y|��{c���_ի��n����'�Q����/(:���x��g�s��~$8���%�ν�������.]�g���Z���ʑ�F�����Q����>_gm����g��_���{k}�K��W˽�=������>W���L_s�ǩ����=���;��,�ձ]X���������]�'6���K���������;W��>�r��P����AG�Yql���<��������/��W�_{���p�ْ�??�v����)�����x"���j���+������ߣ�,����0�gϱ�B=�W��ܘ�,�h�l�����z�G��O���)�oXc���w��x��=���w�������#�?�;���p����u_�8��ϝ�����o���w[,?��,N��@��~��.��h<v,�Q�����u>�	����t=�1Q����G=�d��� ��x0	��`��wZ���uh'��k�#�A}���V�=��z��l��t9�5�S� �f���~�ϓ���8Ζ��2}���;�|~*�W�sCQ�-$p�����n��%���υu^���g�����?�����_��{���T�s������o�Q�\�wU�~��oh6�'���o�~+���N�X�T?`��E����	�q�s�d6������@c��A�����Y󈐷��6�O�O ���!T>d�����;]�c�=�Q�~�����/S�/��u>�|o'�{�v}N}��y6�9~�۲����q�u\�/����Ϯ0�O�����r��{b�_�|м�֪�#?��fy���u��g�'�#~�ѳLp�t�_<��N[��߉���'"���`�7�/����JP_�R6�N�g^OAfœ	�]X�.s�+su>��z >������g�����b+��ﷰ�xy�������(��[����{Q[������v��˭��"8�[1�^B��_��v��Y[�� ����}���}���������
��� ^�q��>к*p�{�կ�y��<8,:o�bm�vl�3�<��_������Lƻ��)�"zt\P2��������n�<��{r~��5Г��o��;�C�ݿ���sW�j�r���y��d�o�n�i���5��+?�~(��򙭛�ό��N��ټ�vY~8/��g�,�*8���=����w�t���^a��N4������F��d��Fߴ_������w�[��x~��g<<O1�p�Ә�H�wo*�w��g
z��{zYr<aN곬 ~�J��������}�{�}�ݿ��D�����|����߫[��9�9Nz��-c�9Ӄ�h]�~=�>����;�)}�W��e�z��8���za���W�p�|S��z��RΫ7���������ꏩ���������~�+����z�%��p_y����_	�Uz7���,o����kr�6��������?�O��w�W?��+���Ǻ�\�3���i�?�q�����������r���߇����|��y�݄����w�����c�}�Џu��;9i���3̺O/�W�w:^:�K;�yL�i��0�}���V���у�.�)�����d����g�3����\~��i�8�ڑ�}�X+�<xA~����_��ȼ_����*�u�Ć�J�D�M6>���/_�s�uK�~~�w��z�l��r���X<M���N������~O��>����m��N��]���?s؆~���<'���c�O��3��7�G��r�n��~"�F�!�?��G�B'�����J��<�t�O���D�{�OX?��}����i�����ΏGp}/�cW=hO�Wx��֤�ҙ�9���~��g9�1�A�1{yP?�׌>|��~����D��z�ی���j��fq�,�;��|�S��|=3��G��*��wϠ������g���m���}L����s�yiЮ꫕��x�<+�O��7zn�O�#�H�Y�P�A�����(�hQ�������<��]��|m�{`�.(���'����	����9>���������e)���gy ��>^���3��s�<.Ylwߠ]�6c��>߈}��u��lN�k��V~Fq^�2������K��sgœ����J��m�o��ZO�E����x�Ħ�J��4����&J'Ǉ7�����x?��a8�������<��=���K��h=\������x��"އB���o�3�c�qu>wy��:1��n�?(���]J�h<��#��O��o�u�9��R<G�A�z������?k�n�Q\��u�3�#�]	!4��h���y`$�`�D0X @`�Er��H�#��1�	�`��������18��=������uv/ݵש�g����߹�N�����U����E����?(GW�U�p�Ln�7��L҇�0���F��Dan��c��Ę?�����}B}������'��/�G5n�~�S#��j'���(S�������w�3R�vT5�Q2���"|�����{�~G�����0׽���i�%r?��-�b{N�{���a�%NͫV��u��3ӧ*;N�>���ǵ>��R������=��������c���'���/���]�s��X�_��Z������u���=c~���_"p�� ��-��@��Ʋ�c���l�LY��T��֏��si������S�k��dz��S/����P������?T~_�7k�NyB�/��<=��7ȶ'��N��ʷS�Ei��W�����U;�OY�*9��d�����S��lspy�0/� p��,��������>|�~��{u|Y���qz����{��Z�<`z�W��ư�������V���!�uv~���~���f�s����#87�b�G�^�?�zk'}�z��i˪y�c�b������,�.��	���忿���7��V�[��^�Or�p���m������Xt��~W?��G?�{��������>�X��S�O�Qԟ�߈X��Vr1�1��mn.b|������t�)�g&�q�{C�����x�~)����c���\�]�+�W��r��|����ğͣ�����\��_�2FI������^��`v,������M�{{t?K�C�������V��3b�\9��ՏQ�ů~�H�;����G��~eo�\.mZ�W�?���su�nWxf8{�34��>���9�����Pz2��UrEǝ�q����Y�l�f�V��4�_�3ȋ�bX_fv����_,�^�ST�v�㭢[��o��/�c�������GB%|X����c�U�����wڧ)�]�n�Ͽ۾�L�����o���#}o�����U���^����B���/sY�{�V�I��p�
����
>Pإ�N�������Scd�Ͱ^~EyP�'���������β�}���gi���V���Ő3��/xu>WKv>����O�r��ٟ�5�����w�S���گ�%�ߦ�Oi�����uʝ^��#x��3Z��b�	����X����ɼu���6T����~?���k��H;���G�WX}�'��Ϗq�X����)�Ǯ�YNg�[��k`���������$�MϿ���{��]�,���!W���E��֞�N��Rj�ԏq]��d�쇓�gz������
�����\������q���#���v��EI}?�B���������o᾽�#bY�~��}�������>ַ�EbLtߓ~�_��:^��� p���Y\}u�����3�֧lވe<N��P8�ȉ���.g��y����>K�����s����#���ӧҿS���j?���=�]��{�|��A���#w�������	۳;r��T:P�n���<���nT������p�� �H�����~CۏD�^P<jgj}�c9�}�t�wx����'��,ħr�tk���{�|�����p��`S?���ٺ��)�T�t��(���w�1-�FaY������`�ߐ������A��O����ϻ��Z�O��+�P�Wy��` ׂ���y��<W`���'��@����Û�x^���:k<R�>���y���/�ř��,���]|�#��Q�/���U>��_�W�ֹ�}�*C�v:\�$;����d����U}��*�Z�����?A�W�
�fQ���jO��a���,�_������\?`̳�Yo'�zF��:g�t�Y�����l�!>־��X���~Mݿ`!Of���/�m��[E�밖��ԼR��W�`38�?��t���n�G?���x��a��)���b���'d�Y�(�e�\Udp�����?���S��i��cЁo*�h{�1�]�*ݔ?3=��@�N�K������/�����h�ơ���qv4j?^6_�}|�F��������1Ϗ<�������^��	\��\�iE+? ��r����{#��=~���Z2��i���Sx��~`��瓜�/�<!Y���}�K�zS���������z���/r}��}ޞʎ��;\�]�����Z*���U{��s=������a��/��{�����G��gE?��[ߜ�+���j����!��}���گ)v��w���wƘ�����Z�[+�V��O�'�J���:(b<^g	L�(ZÏ���(�2����zh��{!x�~�������\�TB��)����w����L�}���U�ƈe����צ���)�N��G*;Vс�e�q���y1%�J�����X�/���L���<���'�����V�|���j�R�G�5O�nOr<*{��'a�
eG�^u>��|���_��|n�>��;�Ք��*o	Ke�gz6k'�rN�{j������s��csK��.�9�Sָ�e߽��׭���*߈Ӂ�w;�p,W��ݽ�����J�K;���*��E�[ũR��~T������W�wz#��g�����\j~�)x��������ٟ��"��&x�k�>�����k����_�C��6�<���p��s����8Ϫ8�y��nj���F�k����w���S��M���R�[G��&�k|
���3��1���H�?�|J�����8�{�>6���ر��?��~�}�ޔ���b~L�s�Ty;��u؛c�o�1(����7-S��������|���=¹�{��<���#w�V�������F�)p=����J���V����G���Y����j�f�7��*{��>��7�iq�K�!*��NrI��51���SjR����7���~)��/�.�|}��7z�D�,�`?i�=�{RT�L�۵��߫񴤛�Kg
|�?['���9�>�N���xN��b��9%�^E��W~��\����Q���y��c{`3�c:�I���n�Sy~�C���?��޲v�����yI{�F?9�W�#�h`ė��}^�����׌��_ԟ��ђ�	�^�c9=�����<���]�gv��iy�����1�桎K�w�8�i>;��o?��2��	���3>c9��x���VtgN���z���3r��4�_�+�je���Q����/����`�����u1�f�s�������/�БjW��q��:�}�x'���v<8������o�~����/J��:8���������t��N��ݔ�
Z2�	��y�q��'�����=	~��Ѣ�j��_�ឯ�Ř!3��!���C������h��	}������忳NT8���#�6���S{;W��T�3��P�Y��юg�O��������=�=��~���󤮶�z���T~!->un;G�!����X/�L��S�@&��+;��=����	�����_���������{n඾ݫ��_�q�_���.�Q8����υ�Q9������*g���	�F��9Y��/����t����U�/߿��:-r=��H���#����(��ve����Ѿ�����ߧI���s�D��n;/�zU\����##�gD�m븵&��j��)��κ�e<��G����������X�G�6̕E��_�e�u�A�(�|Tj/�����w���?_c������Y���8������&M�_��O�+V~ѝ�B�/rc����~�>��|��xmo���>i'���-T?�y�p�i_��v���N���>aC�FҞj_`���j�q.t��{�^������_ͣ��~��qn�eal0����|��¾�|��<*��������4�/�[}�r;k� ����x���v�>C.��g��c���b�)h����3�s�w������'}X��,U���	�Wh��/�����z��G�z�}����S�z�B�l�=#���=���j����3�Y�g�r{��'�/��͢���E�h� ��\�sd~�?*���S���{T;�ڟ���y���T���g�J�������N��*�%������Ǚ�)���7���V�?(����G�_cq�h�q�Ǐ��g;3�卬�(�d|x���������OY�V��sY|�?��н�Wj�e���O7<\w\0Oe�p�\���pţ����wzl����;�8[���A�s\�s��f}���55n����>����������>�i�9G��_�ܨ���)�sN�w|�zo'� ��#HO�c��o�>��a'�T�XS~Y��I����'�a�]�y��؟����ל�X|����/�����;�QUހJ�U�|'{��s-�p�g��B�C�|����|1�_��~�?jy��=^�9��?T8y��F���a/�u1��V>$�,���dq?)� ?�ޛ������%�ՙ�L8|QzΑ��"�~���7���x�i3�3�e���Z-��Ƞ�*�mޟA��'��g�7*y���/���w{��#*ˤ_�jM�H,�nZ�K}��Y�9ק���z����d��z��v��E�m���NT�σ�w[����{3>��r�j��vϤ�gĴ��U�@eoG����nѸ�L�Wr��۽{_O��_���˥���1_���:��ӭy�y�ɘ]�z�¯�O���ڟ�[�=u����>�su�d��r8��,<�	ڝ�� 7l��M�;�p�Ɩ�/���a��y�#�1�C�kڈ弗�����Y���~�����}G�=�s�~�쇩qk���?95��eʹi��o3V��;޿����]�9��>��~N��O���$�}�kf�����H�c��a\?�=����P��c'��B7�N�g��g��_��6�fȱ�s̈́�s�΍|]�|��Ô�P0����jg�+<��V:s��E>߫�o5_��gH}ſY�G9'��� �y-@�����<>sޟ��5���h;i�{�����W�%���a8/��X�?������"�Wu^�����{���<J濊O�4�WD�n�y���V~u�֟�r=~L��9S��]�t;��k��]Tz����w��{{P��1��,��m"���u��?¾B�4��ۊ�h���G�G��܎b�j�:v�sc��{�+�w�'���0�����b���9Ú�U1�'�%��Տ
����'_)p�/��x/t�=�.�����r��C[�����	��?�ϋi���_�iꯣ>�\&�ۇ�ϐ�8���yQ���=>D�������>���w�m��#=/�ｦ?�~�<
���iK�����aOQ��s~�|�/L�6jWSoU�G|Y�:wP���k
�V��1�i�W<�-�q�0j��pݯ���s�|��U���������1�i�W�v��9bY_�oH[������ý�k�}/֎/jMU}��G���~���=���+��=Y�	��5�ϣ��_��;��o3�-��:����������·�������]�|Δx�|S�����yݹ��
<����8�sp����%د��+�<���������?�|��%���1/t��|�O�g���P���&�������;�9�v<;��39���Y<^����h��x�'��x�u���a��1-oy��pQ?�o��|��%����oM��]��������D;a��X�����n�K��||c�g������E;K�U�����~���<��+i�����#�۪_'���S?y|�֯�JO�[̋���~��<���<T�}{=�*�����ُ6Tz/��L���I�o�w�} �P�������}��Wբ�zl�}n,��������������Uތ���\��u��"����B�W������|ɸ��#ې��U�]�$�cW��Gc8�w�˴U|�v����R� *���x�ǱP�Mу������V�+y����鹃Jns/�";�X��ǝ�毿�e��^�����չ!�#Ƥj\�5�O���ʙ�K�;9�$�a�����+�>��`����p����|Yʇ|�f����G4�����?���Y�g{�U�7>_�u�B���=��O�?�sI=nov����{�$�ϒ��ޯ�N=[�������o��$��6�|?7�������gr��l?���=�I�����n���r¿�U�-�;�[�Ř߰fC�/8�}�4��N���_İ��⮝��{���|	�����W%����ywF�������~1-^�����幭�Y���O�a�X���l�i�pm��s��ّ�b\ֵ����2�py�m�#J7�[��~c��;���|����8�Zf_9}�O����!��
d�cy\8���Q���������
>_�|Dlb$u����{/˚�G������$ゎ�خ�u\fW��׋��k��������bǜ�5��ξ�����~ϓ~�տ���bs%����W�b?��|�R��|Ƽyt�)�a���u��b�ϲvj<y懟*���ƛi���'����c�75~���.�{��������f������wM�/iϢ���g���|ڕ�k�Kc���E�'�O�_=/��%�D���8���9�0:�
xU���dq����b0A����ϊ!��||������[�K|��q�?���~i{��ܭ��7�c�-Y��.�rE,�g��à����G�r.�����x�-�_��u+��J�S*�����}����o����z@���O�W������8���;3�����a'M���co�q>.�؆�����{����}�#�C#�O����SO�e}��xg���}��h�:��~�w8���Sb�OP����H�a�ʮ`9��sw'�?�p���8������7��A���u|�6|�o`}�ԇL����eI#���W'�+�/���N�r�4��d���۫{�Ԟg^��[:����m��z�����g�"�֕���2ԟ�+��
y�`W
���ƫ�ۜ�s�-�c�w��U���O4��3��uR&'���g�3��b�O<΍�YN�gu8l�)�Q9�M���G�r��R_������3�ةF�K�Ǳ����>�]����j_f�� ?��@��>�a㽗
���tS���2��۩1ֳG���bqsd�jf�_o?���<k�Y[1�kw0�Sű;~�I�?<�o��y���7�@/������{<�&��5�=1��ּ:�����|{jl���#�_���p?���CVA�k��J?�_=�8%��*~ų!�L��^�^q=[���������+�73�J����.�)����5׫��G<gz�����j�␫���ِ�
����滾�x�#FF㎚,_��@��9Y�����xGy#�(�y�?鯷��T��>`[�2�,G���j�����<����
o��;�1�+=q$?ƛ��8�m����C'���A��aB���A2��w�ܣ���(�/�����������������!i��ޫp�/�������].�T�z�fǁ�ѥ��{��\Oe�8~�gyz}���s���̇��c;|]\����q �xvoϧ���-XϾZ�NS�Ƕ���Y�ޠ��[Wv��:��>��'lZ�I�Gc<���tݪe-����_����~��o2y���`3�H�C�y?���%�d�~alN�����^��YV_�v����Uz�ZT�pw<��w���m<��a����2� �p��w�}���=΍{�r��,?u�����%>����+m����K~��?��V���G���?;�ʲ�Ε]W�O�����k�%ٽTSۣ�7�~��������^�ӟ��g�G���M-5{�!ύ���~�/���1��IǻX��n���_���������6���T~�q�Y;�>����z�{uIR?;D]��\إ�×���l���W�;���w�{_��=����s�7�ʙ��m��c̷�_lx4�W��w8?�}���h�U�y������y����,�{l�uvE���FΟ����������cb��g��&�_i�p_��7~��K�3r�������U1ęA�}K�ޝ��7#}0��~�/�#{����7�����~A9��{9���V��-v��v.�ѽ����Sgv��1����˷*_��c���+��O�ٌ��^yX��?��Y��د3"���X;��U?*s�A��~+����H����l����1��!�S�},�r����E�w�C׽��󚤿������˓��>����|���?�n������1Y�u���	��ʤ��I�Hg���x���g�t8?��[������_�^�G���^�H�S����u��m�������
�	V�	����sK��Y����⸶blW�%8�<�;�L��W���P�.����g���E{��'�k�c9�����:���&�}YR���
���ڗOm&�#���vV��|����Wy�ԞQ<O�gZ}ꯊ�Y��_kMG����J�G�^�{f[s���{��@n�#N�a	�3�w�]#�oN7���P�U?�������gټ���>����ۯy���k<ύ���ð��J���D����%pm�/��Ѥ=�[}�ߢ���������ڣ�7Ǹ�����O�w��Ry���¸d��>^;���]�ž��G��P�\nxX.1��ڥ���}1�?����|���p�����z�p������T�j��V�����1���k'��qr~B�+���фc�v���(���}�U���,�lܧ�u?��x	��|�׃=��5��I�E���|qJ��<r��M�~�<�;�_���+����:����-�}�}��|4�*?�	����xt���9��+�_�a_l������ǘ�&Q</�תtS��C��?�����9k�cc��Ω�`k���7�v,��Ύ����?k?�D���[�_���9y�)�S����A��c��^E�
?�S`�a�T�U���#��������5h}��_��Қ�~�v�|`�^�mU+��7����ʦ�A�����e�^�_j_�=��j���հ�0aw}��+�N\�Řο��[{r|��|��K�#�~��b�\����ϳ�~��6�k��9��� �U~��;|�y�Ϗ��N�Ln(ͳ�p�����f��);=�̮�~�?�_�P���}(yo�ޯ�G;��3�O�d�D�/��1;b|?�X�W���-���ls��M�������Q|���^�G�!������T��Z����&�|�!��a������R�����Tt؉>���[��x�t����t>���xn�ϐ����u���C+?���_��y���.7���	<k��Q8�m���ǰ�~[���O���+p��)���ϼ��R��v�gft8Y���a؀X?�?����u�{�7�����yd��E���O���z8>/���8�}������h�������Y?�ز�����6��Z�'��.'ٞ�������)�3����g���ŚL�?������I��g��|����c�Q�U>�~�W{���8�Q������+�役����K>�yG����Cv�|'�����A��)���߇=��GGb�O�v����/���y������=5�<K��^�G��F·;G�WQ��x&�K�x���c_u�"b̟��]E�rrx%ϣ�󖵇��h|��W�{Ɵ>߫<��K�l�|]��?/��1�Z?��\�q9\�ޔ��:�?b,籮~N�*^�㕬wf��Ñ󏮧>��C��_�>�K�Wr���Qv�����z
���~BR�6��#������ǫ}ƭ��������cꗮ�ר�Џ)��(|�]���:^�;������|	����sy�q��������,.e�|:V�^����S��:���`l��'�!���u�O۟���/�K�;4ޒ���횷�~v�!��c�G9����v�o�ų�������yz���/� ��L�:�<�m~K,�k���g[�>S�N13��ܤ>������w8䛮�T��<!}N��}K����_S�A��%�h\�	=r4�ϲ�n�.��&�|��	��?�ϯ�Z�dr���\gy�=��)��;���c,��gĞ�蓌>�s�G��)�{1�?�����K�3����ag�������ε��S����Y?帝Xksm�����v��Z��nߒ��o�vd�V���Uq�պ���*}���~���Χ�����ڏ�~1ݍ1�;+��L�Z���ȇ��J�j�w�Wy���#���x6���S�����+μ�g�Xγ8~�<���}:�u��z\Q��������Ƌ��O�N�,����?G���(�qT��c�X��|����?����"��9���_�9��r�z>E��O4T�/|OC��������yB����w��1�L�/ rZ�#���˓~�bY�<��1�+p�t��:`�H�L�w�xo�����,��������b��]�m�����wE��n�<��1�U�����?���x\*To��{⮏<O���v��<�?�o�%�'U}���W�kc-���G
<���_
|�����/���y�*��u��ñ-��8��JO_�0ϫ���Ѹ�y��j����q�}W@_�����Y��>�ñ��4<7���~�z������/��~o��1�c����[,� \�����E39�~�����#�y.ՃS���i,S���NS��[Ovή�+��)��oK������ö��N�/A�~�>�gD>_@�CI��������a��n�1
8Ծ���=A�/�]�W����M�W#���~C8ϱ8�V�o��]E7o�E����<xu/��9�ـ�ߟ�WW)�h��%x\U����7�w�X�^�k�QǓ���Ƌ�����x��?ޟ��y�c�Q��l�_��0F�q��'7	vxz�ñLO�֒�O���9��ݧn�7>�X�����N�8b�s�~��9!ߞ��AQ=������c�j+��M���ώ�]�4P�T���*�q�v8qU~�'�������y�����6ϝ8�D8�H��G�����^�?x�5ĸ�������q�����'I;�R�L:{�����ϕ>���鿷??8r�������{x�~c�s�jϪ�i���zh'<�,;�G��P��a��u=��4������Qx�O��)��b�%Gc|~����[Wu����#��o���cxm,�jYI7��G��c|.@�q�]�X�G����rz�����u����}(�?Q<�˜�Y~�jݟ���������z��W���Wt8����،�^c��;�M8��Ü��*��β�����b��z�=�վ��7Y��=�Mߩ���q�c�AYE�j��T�f�~��[��>)�����|u��1 v���w~X,��1�̚�_�+��W��S�-�������;zۯ����|��mx~������Hy�5E;]�����L3޵��}\Ήm{![9��K�8?[���F��ugƇ��[��>�6��_�x	mgF�� �΋U����!��>Q�=j����4�y�δ��}+�ף|v;g��o����~�����C�ȁ�O�����C�O����#.�/�ϰO�|Y���v��c8�/�'"�utΚ��h��b�����,��N|�p��5NX�29��F�G��]�����V�31�25�A\�K���s�׻K��}^�1���:���kȥ�� ��J�c�;�%�~����_�~������aJ}�&�m̋��2��6��_k�$����X/hu�3��?F��yG^ȍ�n�������ց����ƍo$��=���c9yH��W�5է�u�#���Z�w��1��� �/���,��{��Gے��������Kc,��w`'��}������;�c�#u�^жL���~ޣ�z��_E}�S�d���iD�
��S���y�ho#���s��Q?FD�7��վX'��Ol��?I:(�I{�KR�����~�����ư���D,.g��,>����I�L�1�7��3�vf��U�������o��u�1���������?�����	-�\S���*�3��u�8)���r;�1�y+���j���i�_T����W�m՞L/ �[��?��Tz��{��F�4��*����|��!w����vŁߌ\�����Bޓ��VX������.�������:��+���LeqS�����z`o�V��v��������>�_�s>a>����?'bX�AN�<�x���GmU�{��u�Ù?�����/��t}T�y��g��3������g�l�]���[��;�v��m���o�t�#��ۼ�t8�����q�s�9��O�u�5_)�u�-1���q���:������;|�~$����~!�O��IX�a��[o��6p���T��j}�����3ڠ����7�y�0<\��3xE�����u��������;����-�}��)�g󺢳��1�k6ou�n�g*\�m���N�Ǔs��qS? l�a�����/wŘ�#����b�7o�ۭZ�����[�*ic�NA���9�V���{�_��:�g��=��>�3���k�U�K��L~IF��#Z�����EZ���K��Ъb��������'¹�����m6���b�nn��������H��e�a?����)�O���V��f,���k_�w�e��=*y/KƟU���_�WAo݇:����{��-�ńS�����+���o��VwM��{�;�Dn�f��:�3��G'�}�x�sg�Y�)����n��q���N�ݲ|�.n�u�^V����<-���O��~<̹��?\����{�U�~�'J�*��G�[�y��A΋�N�<i�t;Wp9~�[.��g�Xނ/���ON|�����w���uG��V����ֹN����Z������r�W��ѽ��u��m|Y�{C���=;�}U�T����3w�8^c{��'��g�>��}e:1����c]�or�?g�;�C�����������4�Z�^O����&��>l�S�clo�:��_�~��;��y�}p�ՃU�*��α�L=���+�G��n]����U^nk���wq��u��W�~��v���GR9�������3��%*�3�ӟ|�둪����?�Y�u���r�;i+����
r���������vVtc[WٟZ�����������C�]����|�h������:%O��iY��f��e!MԮ8�?��o硟�к��J~�ra�?��SG�q�Ġ�`S+�V�U�N9�����W�B��~hk�5���5�+#���h ��~W+�_X�!�]�r���q[E�6�yAq����V�rM��3=����
g�]1���C*vά���Gb|��S{ݣ1M�c{ͧvԪuh��v�/S��w.������o�[����Q����woƈ��";����X�ٞ)ү��-�Î����}2:�=z�ս`��x=��1�{�\�{$ig����~	��zML�{��}���~�*���gb>j܋����y�ܧ�<�jO*��Hĭ����i��|�`������}�J�W���������,������sH������=\����2?{�������޷[clǞ��/�}�w���qq�h[�u��ЉW��;��O����b��s�q�4���Ἠ�^�r�uϣc?Ӿ�{���^��
<g��	C�۱���O:���.�V?6�yh�d��a��|ev��uW�ޫ��֧����������nsd�W�x>�?�uz�J\�����8�˻N=25���~���W���K�#�n�q���O)���,�o:�/��JΨ��������sU������ta?���h}- �u�u�ñ�<���~��v����������R�:�x�u��/�>�7����N6�got=U��X|]�qM:���I�n��vxoƶ�{=>��{��s�M�����?��j_����N�{4�u��3�w��1�����iWx|B[��=�5�E����|��~��a������~�T�]η������@���������ۜ^��A,�1��#�:pc�!}2�Q��Zw�'�~fؠ�<1i�Ny,3�֙Q�3�x6
8��gF}�_�5�`f��d�J�������������C�V<����v<�ߟa[d~ݪ_.?�nu���p���tPy���w��ҟc�yD�_l���?���WM���B����i�꾡�*���#���}W�����ֳ���ݨk�U��R�_7���~
�sŇ�Ge<m�U�Y�_�*���ɪ~�XnT�1o�GE�@�/��f�3.7V�-��w<����t�rYF�*�N�������{�gճ����Ϡ���J��z�J��M�Ϛ�8����T�{�Կ-�u2��3byܭ=k�����g���|��l��%X||/��޷���I�o�Ӝ>��¯�r�������+�u����L���D{�O�k����ǐ�t�>RX��=1�O������q6��|����N\��#���m���,S��l �@?�>�,���ߋrVg���0u?����a�"��U1Ϋ����/��A'd�{���zA�0w�8��	�ga��U���k��G�~	�3����;�?����}�s��󨬚_S�C>�uqE���>��c@8�B���C|���{�Wj�q#���g�gع�"p�{�z�m�� ?W���I�y������ڬ�^ߟ�zz_�@���v��k��W����������$���{�ٻNY��?�_7�t��fGU�����9̃t�X������sU�G�wv�Cj{*�����ΕU��W�4��`ٌe���G���Η��3�c"��>Q����Y\�����п��ԏ�כޯJ����'�;<��j��֧=��1ȋ[c��u���<����/��K}s��Y�Y�/uxe�P�O�}���W�wS�Ɲ�+�j
����M�N���v�o-���C��y @��btO���V��἟�:��k�YÙ�F��F��_N�[�K=!�V��>���ә�̾�����gG��3<�0�y�.����8�ϗZ�*;�¿���+�U�y_oR��8��:�*�ӏZ�Oy�+?��Y�9��<ȿ���;bl��X�q�'T��^�	����$���s�?��Y�W��{D�ᎄ�&�u<���1�����!};v����m��Y*?pE�O9R��^_�{�g2~v9V�1�`�ݐ��	G�D���%p��sy����ک��}��pv9�5��%=��%�����Wͧ�x��H_��|s���1>�]yyo������Ķ���*�H�{ś:���|)���������u�Ǔ�<�������ϐ-�A1_�M�^�}�c����	o?��������m�|�z�,�˞��7c���18�T�]�V��X*�����=��n��\�O�a>��v�h�i����;���G¸ 7�ת��_U<���:��G~3e]�J_�W��b�u=��Q��[��(��x{\y��ۜ������.H[�K�=�C��.�?��_�<�q|v�O O~)�϶fv��i2d��|���'w�v�.�`�ԟ� �i������=;��t�~���y��^oW�r���O9/���O����C&��<�%���	�i��ua޳KO�_1�{����p�7*��r��spw5<��+��z�,_����0���9`p�S���{3}���8���������<�ð�Z�;���X�;�^���*�Wߢ����}gU�U���j���{#��F�Nη�x�C�Ǭ�C��=���W���Z�����c�����Pү*^��G?�>�|F�loR��Xŗ��ќ�'"��2<;���@����.张�(ӏ�/�\;z�_�W�����[�ȇ���U;i�P���D�<~�ݲS���W�u�����z����]�g���u�;cȯ�3C?.�o�a�!f�<��&������k����/��S{��:o?��A�&��H���:���st}X|���x�����kN�L(���ծ;Y>d?��%.���Ty�3�Ο���uƫ<?��T�s<�=m����a�w]1t_����gc�얝�d猲u�,����������s���꽰�p�vݍ��o�_�#���>#�B�;���1���݉�?n�!�O~���T�8�2͇�mT<'��������V�����e����Ͻb���xD���w�y2��y�U�%W�?ܟ�:��w��~j��Q��3ȯ��WL�w.��~��ծ@޷/���Կ�Rљ}V;���Or�K8�.a����y��П��0�4.�ź�K��<�	���J��N�G,�/m��^r�����ۯ㾧���>��W�.֒��J�:��O���߇��G��p嗮�C��q�|���u᣹2�/i��r����|���I�}֯c���㧴Q�����5��Ø�=S�9�[�s=}Zcx��,�ϧ\����j�z!�g_'��:n�~�����52���׭�}�8��r��J�q{z�*O]��Aq?�Vl����uY�J/�����c�.q�9����9	~������G�G�_�v2��>Q��)� Ke/���N�8}*;��`���/�'T�� ��ݐ����x�>��ok������|t���?:;��*���O]/������/�?�u�W��`�y4�_��~`��7ru���~kjo���t~��u�f~��1��S'�����ո�������z\���˾ی�:�z/l[���8���7��������{5�5�=�_����~H�k]��Ur��_�O��{�U�b'+2�5�y+����#6	��0��J�{��c�q!���y�t����GyG,�<1�6�V�N8d��N�/���Vq�S�|-�g�[���R������;��T��Ϋz=�²�ĩ���ϫ�F���V�d�O^�aXOe�݄���u�:۹��ϥ=�_��u|�������>"�O���?<4���Cs��t?��պ��ϗ�g���k�'j���3;��.�g�(r~s��賸C1o�e:W�nѸ�U� �wz�/ߝ����'�^�_��(��?�`�{]�~��u�+���1��b�����#�w�w~Y��Iv�yx��_���z��w?����x�p�^�'w�B������kc��x,���:M��_`�0r>���}d�ʏZ�w��)z-�WvȪ����?�}H=7J�\�]Tq�_�9(x)���~y�Ov]�g��z��¹ϽY�O�Sְ�p��*=���x^����V�Co�I{2������ι��˒���<b���~
�0ස����b��@�9;����u�±�|zo�W$x���]���8O��u�b,'����_o��p#����iB5������{����j{o�Syp���y$���A=�à��s�Z�����v����������'����ڍy���>8�wZ��
�֧_��1�W�u\��|>��l���*{r�b8t��iO�I��E?/�J����|G�����������R��^�v���|������b�����,�������3����v?�~?��{�>���w���`�G���m�,�5�_���/��W�1?m�W�We?/0<}��ۂ���X{�o�|�=/�Q1��؆�������)�b�;��֯#E����Q8�B�������8����1���%t������e*oC�i}�����K�_������%���*�N����h��ў,�9"�{������~J���S��\W�g��yb���t����O�x�PpV����k׆�C�5�^�r���;Οչ`���}���_�G�7��L��{�A�l��l?�����	~���>��W~`{�X�*�Ӕ�N�����{<r��a�����ޤ�ax8������F�Y�/��7��}��z/R�g��:��Jz}�a�gn�r�������~�����=p4���@���˟*����f���L��t{�����3��2������g�/�y���M�?��>�>���2x.p��}�]�;�,�NV�ef�e}�Uq �z���B7���̐��}���S��Ͽn�; ��t����{Y;��k\P������Wٽ{�E�>a����yg,�K�rR�<�?_c��4����錹 yY��9�[���|���O8��W��'Q��l���~�����1�Oc/�kb���8�N�|�|����i���;���ҿ�����������F,�������>l���Mh��������V�Ռ���oQ�Jg���(�+��\�C#=����>O�)ϙ���S��O���A�*�Z�w!b���%��=l��9WqV���p�J�<������_�1�O�S�G�~��`�|�v��]�ou���c�w���vV����H~c��UvȪ|}.�����h��r����p���N�#�v��cl�Tv�E�o���n���d���7F�ټ6����?�Y�N�sd�s�����_���*�y��;��O��UE�~���}ү0<|�����ˇ���a_G��~~s��C�U/L�o���eأ�|���M�'�����_9�7��N�*��<�����h��9���jg%��yT�mp��˷S^��]:.��z�)���m~���ԧ��<�o��}�O5�L>U�s���������2�ҡ�?H��kz=�S���iG�/t��_���b��GcL��sԮVyX�7���9��z��1~�e�{���Ʋ���L�s�>�����ԏZ��4Ϊ�7��O�������r���ƚ��cj��O+��G��w3�����S�x����km�v|���~�'y�N�X�b�}]oVt ~�N��J^Uq�<a!��I�N�?��Y%����:@��_y�����չ�cE�.�W���>��*���WH�3<}*y�i�U��*���O����xJ�S��y��d��1^wؽ��&U+�]��`R�}p��m�c��9����;�x�?���]�!S����,��������xc��oV���;��+_��}O{��?��1|Ы�M�Yţ�n��]���X�]���}������.����y@#�ÏEN�Jj;!�����^���6֔<H,S�Z2�bH;���:�X�ߒ��|�8��U�󛯧V��}#�C.W�;���:�{ë�s[���_B�?��g����B~>c����#���1����*>�ڿ
���]n�ϐ�g���7��{���󤙼u��<��~w�3�y�v/����_�Y�����+>��_�ʎu:�>�J�8C���*���b�c�����	\���T����~[����|�;�X��q�X�c�����'ę�L��#��l����#����{OV�YG�_��X�����g�����n��/����k�(�/Z�3�sC�}:�ly���=�cC~��n�{����}�}�q}�NQ���r(�x�꾤j|�uGe�;���\�-�����*���3lCݯ����ן�ሱ{kҞ�e�����a���}���*���l�u��&;��t&W���'�����Ż!�'��?�|o�GK������;�V���;��k��ǚ�P�ح�q��t9���Q痞C�������G�_����1��J��{����۽:�_����
��}zl�=)��]�w��{V��2�N����C�мI��p��V���;���Χ;}~�?���OG�N�C�Y,��1�G!���?�q�����f�9�T�����9�2~���P���u}V��A�%�7Zfψ�]:��]�w��f>h�j\���)�E�K�S��;*=�%���H.���`�Ή�'x<~����3�S�]Z��7��z��������;4�+���3�?�T����D���9�,?I��j�����ڿVݿ�������w�+T�p��S��,;�R9�5N[�,����W���z���IS�O��~E]�*�*O��K��g�1�K ������]?�N�K�[�5:O�Z>����?W�g���z
���z��cR�g��|��/��{�����B���I���	;?W�xY�w<��|�9؟�6<���oPK6�'�O��V퇜D�"���x������W�N����|�v ^���U�h��ݟ1��N?��b�zE�^���z������Ǳ�=�O����弣��i1m_��[��$>��ò|η/��.ȭ7%�}�{<��Bܙ�?+=������<��z=̙kV�c^T�P�?[�����V�]Us��x��Ǹn��|=������iyVW�KN=/��������*{��[��/�8>����b���=;ry��mz�@s��}�N���t]��/����^������s i��1�>ḓ1��[�l�@���ۛ��{�Z�gh˗��jx�K��n�v�M�?���Ϗ<Ou�g?�����üj�3S;��_>�g�r0d�U�W����8(�n��mS�Q~��@��y�zA�YS�gt���y�ZYN�OX�[�����N_�>��~3��d�w��*{F���U}7u��rw�?<�%��=ܧ���%��y|Ku�B�������g��*>a�~P��(㾸��S������c&��?�dX����{+~�*�V�v�7�ۺ_��aQ��b���ϩ�����s�1|���.��~��J{��G~�,��FH�;'���t;��d~���Y�����,j�d���y���>l'�9`�j}}a��nV_�^�>�dgp��H������W٥�n�w'_tJ,�m��>������Ǻ��|_L��y���,֯��3o��ڭ�7�O�/c��]e����)z�q���O�	>��Q�������S`/k|�N�E�8p�wS{)��S�@�l���ۮz��{=���O��Ϲ�-��e�	I����^��V}�c�����������q���-����q�\���<iǄ�g
\煮_�g��П?i�8����r6d��=��<x�Y\n��a������.U}�w�Wv�֧��>g�e�����o���W;m�|���M�of��w�"���U[�_�����м*�������D1�w�ݭ�?��mv��3��*����p^x;�c������/�8O�'"�k���z�.�}��e����O�zn�T�'j/e��x��;�_&���1��ƹ�}I���kS�"������U�}�}�/��~ ~���o�3���#����8n���gŘn���N��]���y{��[�J�?�홺���/�a���=�g��K�������,>O�v�;�ͮ�G;�qy��$��;=��p�+���VҞ��?þ[կ
m���c����}�����=�����~!r~���%�k���g�yC�k�����1I}�R��t�s���s(z�R��t8�W����~q~U�G>.�U���������K���m�uD��P<�;�P}G:x�vw�{����c��oM޻��������5�ȳ�߫�8_��~��֞�V�+���Uzv����:��/��|_��^�?�W�e��� x�nI����Ws���o�}�sk��F�~�cx^ٟ���#p���1��p߿��(����@d�0w�s��=�3�\���������%�)�qތ�Co��d��*N��ر����?���	�W�V�E���M�m�����U��뙾�;��q�cL����~k?��>��N�[���o�|R�}�#�w��N��/������ĥ��~���y�N�O����T}�~�,O��ܣU��X��X{��G�NP>�~9|���V�qo��� �ͮ�>�J��{^��R~5Zz~�>�������V���6�6:l��Cg�Q:?P��5��1��o��MX/�kD^S�����y������w���?�	~�+�71������������Z�_k�%�EQ���g��f'M2��a��C1�4�y�t��*^��x�ٯӋvVv����^���=�yr��������^��j?"�۾~��#b�.���8c��x0�?��qM�ά_;�c�qwj��7N7�?�='��y��ʟ�t��Ku�0�קY;��}��}���������V�w��i��sf�O��5{x۹͗�''�6���]!�[z�.���ݟ/�ϫ��˓U�1ϣz۱/t��2<nw��fu�E�0>g��9�u���ռ�u7�ڥ�f>�	��a�7��wW�M�XN�k��I����󛨏�:9��O�~�|�|��8�U�����w�˚�]�hQ?������^��K?˦��ȼ��2<��9�1��;��8꾆�-�~�En�^8��Ӛ͸��S��yƅ���=apw�<"p��ҿ�sӕ<Ḻ?m��^��|_����LV�V��c��+�����Ҹ�jZ�C��W�g���K�����_��z�D����rg`h���̿���~"o��O'�#[��������o/�e~��xs|�������gDn7�28���?��'����!����b}�M����x����iQ������xib��վ��Y{��?h��E,������*~ ��V�1���f���U>�����U}��]Q����c�^������ϴ�<�Q�7?�j�jU����#\�ϟ�C�gv�����B��ҁz����Vz��O`3��L^y\4�[���/�x㊯��y'�O���xX6�ϙ��2���¯��{M�����-�$�r�m>�=a����A�ӏ�v��W��9�0/�#pȜ��Ӹ/��O��5��_��S%�>"M����4y��|�l�<_�����=��S�?��_��[��wů��j�P�G�|�g�*��<��p�Ϩ��*y�%�72��|��=���1>G����<�������V�g'�T�晜�b��i�N�u�V�G�����~�U�=|���W�?�Ol�Y��׷��!J�9�U��Pǋv�О��+���Y�Σ1�n�w��q�|�)������+��/���=�Y�S3�-�3�G�xB�w�s|_~���#y�<on�kb��i�D�{+~�Ӹ0���z_�%����
�ۺ:��Q`�e�[�S��+�w���c����u�y��j}Wŝ�݄s�>��?�?�?��߹���N��e1��T�W��r=\�ݹ~d=���/��r9����V󽲓7
�� ��;ڇ��gm���������N�Ә_�%�ݞ��??���?���3�d��S��S����j�����v�����_ٟ�y�{�>e�B���@z���;�{������w��!�wN����<��-?�9�r�sgn�)��Y���M�\Y��)�_�.[��y��~�=��<�O\=3�S��t�;䪤�����=I�]Qߗ�чs9ó�x*9S�q��*�E�{�#���:�v0y�ϋj��}z�{��x��<��_�@���L�������t�Y�+{��������p�ߨ�pX�>����Y�<��%N�{:U.Q�W��������Ӈ�>x�6mc$p�W%�+x����s �t���"�美c��2��7<��|������L���vk��R_��}H9��yU��_�ͪqQ�����ֱ���{+~��v�O:�}�k�*�G�Vz|�:��^ɇj~=$�����)i�Ӂ��A�O��2Q�|�J9�y0��b����U^�c�����ֆ�c{wG�_����������'�a�o�=��N��o�w�3����v�/ο����� {E��#/gr���W��Zg�����̰��R�ï�s
�����?�6�������cؿ<��������@j/���ey�y}q ��qjQ���c�x���r�QI}��3�g��k��2��%�c��]D�^ϧQ����u]3��K;�㇕�~���[�C�FYG�����G��������<���v,���18��c#�[�S������+���a2;��oa����j�5S�c��@��Q����O�����/]Gdt��L����;�c����\ݏV�oW����_*����<��{�C��-�c��B�W~$��^�;�_����*�sV�zl����ؖ!'�g�yT�;��>U�$��[��M~�����Wb�yk�
�h�w �����c,���p�=9������'��ڟ)�:��=_�_*}�_�s?W�y���#��~�=��h���Z�y���U��ǜ77%�����	Z_�-d�߭�NzY���_�y�9�B��yd�s�w�/y��/�>K蜧�2������İ����v��Pz���e=����vc��?+j{��K8<W�P�:���W���!ׅ�֒��gU��{;�FA��V�0�o��/�/��f�u��1�Q����������c�\����������U�W���S�/�i�����֧��|�s����S�Ő��~jL�*�����3r�a̳|�U�����{���|��W���oߥ�U����c=򼤾�G���U��:�z^F�4GfE�)� ��U���>_�x0w�#�/��^��ͣ��+��|��X/���v0u�*>��w.��V����}��|g��W�p'4��Y�����0j���D|'_��A�����S����w�'k�5�K���@��-p�[lZ�����~�O�ɱ���s"�#.����Ƕ��5��ey�"�|��8/��T�	�m]%7*:���aC���S����7�?=g�mQ<�sl�����a�Mg'
<��c<#;<Ӄ.�xκ��N���1��k�_h�V�g����~����?��٨�����K��c��;<�e��?�0ȏ*���i�b�얟8�2�m�c�q��u��~��ݣ�턮<�ͨ~�� W��� G3,��w_��]������ψ�V�z�^�cy�q,]�,�Y��;���8?h����ي1=���1nz.���{�G���зu��g����_�����R�c~>��U���?��KT��'Őt�y�~���xƞ���W�c��.z�n��ǟ��?7���%�t�<��(ҏ����?�g�ׯ�X��Q��se�U�����N�Ƴz{���ڻ���h{e[3m�y(⺸��v#�������K+��3�J����1<C��q� �d��]��u�_e�Ƙ��\ڍ�����w8����לl��=��R����c/�u�y1��5��'7�7��Ξ���j�U~�G��GƤ�3�|�����h���yD��^rC��}�yG9?x�E��Τ�p�Aq+\�3��Vvi�`F�5��w�L�3ܟ����>Y�v%�����O��������f���q�����/�������Mڃ�ꧢ��ٚ�/�o/���������l�U�A��V�����n�u��x��c�o2����l�;���/:|������vx(���o2�4ş��z�c)1�Y���Y�����L�[�/�9�<<?�&[M���*��߼��!����Y��:|����ǯV�U?V�p�[��c�;�����/���e'?���c���yţ�����Ű��*]�������?O�+������~�Oł�3�i\n����n����~�uM��r�G8l(��1n�1�E�����M�.r���B�u�Q������|\>Qo_,���0a�f�����`q.�ǋs�pă�����|������'}/�C����cp~W�K:�z��w{�ס��΂�M�U��{������Bv�Hڿ�?��b�����ٽ:�U>ï��Z�9/�����{����c���I���s�_�/�l��3�U~�w;�+e���	�����Y�k~]��3��a�O�s�Ö���s1�P ���T}��d�ȱ���>1^oV��tع׺
���~^���%�~�c/�p��o��{=ؿ�ya�~�'�.`~9�L��O��o+����{�r�{J�q�<��;��1�G�7yQl���_�#9����s^ټ�:8��
�֕�����#�|_S֧�3w������9mL��{6�:��mz�S�7{e�q���q�}�~~��FyR������;�i��z@��/�}���xh?�oU.�<�������x��Gb��(����1}.�e;�jO�.�pOv?�pW�^ݯ;J�~�H�SwM��l��1�O��z��w����yC,�[�7��Ý?���~�S�C~��!���7[`ϐ��_����τ��+b����P�G��ƸM�_n��lE�'t~���'�^V�^V��ב�Cw��3��s�{UyVX~<��`~d�2չ	����N~��Pk��F2��zQ����X��0?���ɕ|.��(7�'Q��}z�bL7�+y��[��J�3�8�T��:��~�?�vݝ?�	s�B�{�C��7�x����DҥZ�Vq��̎�w�4<��ߡX��>by��ڟ�������c��|�I�+
x������	���ĕٟj���}~C�D�2i��{�Sս�;��H�g�n'<���c��	�|���l��Y�U�������,.o�?>W��=���t8ڟ1���}�������Ų�[Ϸj}��]���_����x{�O�b���j���T�:�a��x�rW����q{�����
z��[��*<����������<zs�c��_��m����1��:�*}��y����{�'�Wr����ϊ��ս ��<�y�{hp�M�~{t;b��\!��@'7�hv��u_[۩��U���g�x^����� ������|s��'৷� �D���m*5[�?l&�����K"_��{1.Ͷ����V_���/�#@g�︻a�X,��g�$t`�V�c��Wx*;|1�ބ�=�/W޻�����q2���M��9�}:xo�Ϯ��w�b�n�_ǧ��o~?���۰����1��_��hO֯��������f�zI��g��y]�ez��K�k��*W��L�d���ͩ�:#�_���\�U��~De'k��Ӯ�����D.'+�T���X3=0�_�'�~�9��������S�*��"�Y|^�?F������f����z���S��Ca��ud��s�2E?~[l��t}��}I}-�|��.׋�j7h���� ���	��zP��4]��'����s���ϻc�~�� ��b^ �oZ�E��¯n�כ~�!i�������?D��z�_�����.%�+?-t΁�n�r]s���h��Ž	k_"p�y��{�/6CBđ�QgZ��d������/ ��K^������/}ܸ�3����^���T�W���m�_�����fC�]�O�Wz��zM։3�C�y|���:qo��V,󏟳xi���c|��H2梁��u��ǘ|,�����+S�p>��<Пy�����;*�3u�c���Xo=�|Yw+޻Sރ�O>E/Wq�,���o�o.�W�f`^�w��h��소�yQ�Kg�����ž��_�����ۻb�#�o��:^����3��]�휁o ���i��|�^���w-�Pͻ3�~��ABi��ꩌ�qq��/_���5�L}�É�R��������W{C��Z�n$p�ﴹ�R�q>��y���u���#��ո\��g΍�}�|g�n�䳏We�.����*��������Q����.u�;�gW8�@��>�_�`�Ǘv�FL�;|������T��������'�������:�JO�gSzr|�bx
>Y�1�n�p�	Ԯ@/_R�W��8*�ɯ�gFK�w�nJ����Sc�~�����s2��<��h���j�����z9�/������Mϯ1n��O���*���d���W�`�v����7�'���p�Ʌ�ݯY���?����$�+�������H���M�+����ǆ{�;T_`��!�t�^���Z^{Lo��u!�3����x.\�I���'����y�|�8��{��tï�����u~��w	�@�d���P���e�J�O��הɄ��˝����bƽJ��,�����r�e�|T�e��.ou��x(O��OK�{��/��So��tmf�U���UN��
D��스�>��q��L�_�����sX����������2e��=��O���oN��dVqs�s~�O�~�,�:�����������3�|�7���ߊAF����o��G���?����D�lgruqOm[3���䷙A�~���u��i	~�S��j7�r��:� �$�������W�8'�cy�xw�C�9�[F�)֤��sqZ���k��5���dV�a�O����<[��7<�ׇ��U�H�9+F�k��1�e�v���U�+8��y����oy��փ�:����� m���gh�L���>����K�R����u�~������\e?L��<�����I{����{�~���~����~}�>����a�g�q���ϙ>U{cU��5ᘃ����%x�*��	�{�>��փ�yw�dx�}��=���1M�,�G�����߱���Wo�gQ�L�=ȣ�l��O�ܟ���7�nZ�����GU�.+���u�g~��[��;�\��`m��i+�u�<��=g����^�?��*?���a{�>.g>�?ï�����Ani��U�7�����X�Tvi��Y0W��O�
��PR�����:i-��/�\:ߒ_7���~�N�y�)�G�?۟1.�}:�o��?�9��g~ ?�xc�_m��|ګ�*�g\�Cex�����}�7x�/u<����vfy�Q2?��1^����BWg�H��k�����7�g��J��i���uze'�=Y{��Q�s����G�߇b����*?<}'��N�w�Q}=xFg�_ٟ�Z��������%����h^G�8<0pc�
�|i���K�'M��;~�k8���by\\����g���rR�d*y��|�<���ӓ�(SΑ��;|���c�~�<&�ב�x�����~�����|y{*9��>�hB���ϯ�q>O���C�ɮ38��kw���L��q���?#��3�c{ݨ�:�s"��}�������솪�ɍ��X�p,�s.��J��y�����e^��S�����y�lE�	�n��X��ǱP~���Ǩگ�E��?ob��[���$��w0.��4~[큛c���Ʋ�
���!� �17��@8�q���M��>O�/(����~������y|�g���WD~De�9��dg�b���H�����O�����7Nh��i�����s�C���#��A�_J�y��Ϡv�y�om~�y`��Ϣ��~`Č}F���ă�>��j����^��ٿ�@�� �R�_�����簅��nP�#�!��/��l5�'|�\��8����=o����\ρ����C�_�87����+�҆U����E~��@��+Zիb�/1�,�	���>�q�x�g�_��_]�������y�_�`. ��҇x_ext��{u�/�i�~g|�F=�o��W�2:�=�G�"����:/>s��{��R�3"-�oI#�37v��Kyu�ޫ%�>�9�/�������Ƶ����M1�×��czr���Y�<5���u�+l�[���qu�_�?����3�w��������`��k�����h���o��*���B�,�<�������i���)�.�ܘP��cC?f�*�׷Wbo��8{������U8��qP���H��K�u�Z�3�5ⓩ�!���0�Ox�vr柜E�gx=����1ț�8x�;��|���t��C{|M�k6�ƉX�����K
o�#�D��`_�&��e	�j�����^�c�Sl���ڼ�Ǟ�އE\�_���c���I���ٵϼ��H�׃���n�q^}�O���u��5.V��N���;����+���q��Z�j>j�a{*;���(�??��E��ƥE��{~9�s���X�_֟=����c�OO����ʏ��m�{��jm����)�����`�V�F*�?� �C�9�~8���Js��c|����(S�+<��v���_�X���9�\��d�;ՏX��N���U��X�U痫��_�?�a��{����@�֟=��*��w�b;����ZP��!�3C|��/����?t�ɰ��󰨣wKp>�g8?��R��W�����d����s���[&��G0��f�����Ch?|טw���"��K�=�����'�s·�ό[r<�c��'��q9��@�J�ɬ���_��oi��8(=ϥ��"�����m����g{���C={E��M����������|���׼{��(='��Q�'�ψ��y�u��?����ۊyy��+���C;���p�{~>���e~�)�'ӿ���8����=x^���4^��)c���s��ؗ�$��,���;�ͤ��wVvNeo�� ������G�X������bb}��p�H�;����޴��}���ոg���mA�=d[&��֫��+�x����Lh��'�;>������a����k�wX����-1�t��t rd�K��G�_���9�*n����hm�5Y��Y	�ݟSzҿ�~B-ټ�C��v]eO���]�/�|.'?��c?0��y�.�︓���_J��_���G;h�i7R�9��ϩ��vr9���{]��1ryR�w��}���e�m��
[��X�ù��ڏ�2"��Y�ϥ�o�4�Z��C������4��!�s5�?�~*�K�g��������?��ۣ1�W诛~��wJ�U>g~'�eK�X{}8���_�t~��'���>��������� �=�K�?���}C;#p���~��^�(�O@�A/]o����Y������/���YIO�(�\�j����[_�]�uG��~��ͭ=��u����wĿblNİ���{�/�������S�bI�q���t�}z�w �S����9�{~o���p���x�i�~��ZW�<)��l4v����?�>o�1ߞ�7�|Mu.����8�����mzq�gb�wy�����g��h7>��I���u7��S���q���/��u7��W������������k}�������Z�����@o�/���?�s�p��?��,n��;�����/E���^�[4�D�n�|����!�x��޿L���O{���)u?9����{c;O�����W듎�D��E���j����z��u1��:.��k�j��6�]�y:g��Vviu���s<�c�O��/?�U����S�*WU������|����;�����e�������W�~�?c\�������9�����7;�����T��;��6�ҙ��`�O���#p�����E���CN���N�Ӯ�Urc���
�u����:8��Y��΀C�������b�>��W�x�]��
�м�6���	<��k1��v��q?L�ǀ��6/�'��yQ�^׃M�~;�з��T��*�\�s�X?�n-��5E��q�`̳�^���<�����<�9[�������_�P��VC��
�{=�}��M�C?�#��xv���\����;�|�^�Y�֩~��p>�:W��T~�����C��eb
t�1�3���?�69��g[W�Oe?�8�c��@�#�x�@��q�{Q%��܎b��1�����&p�K���ǽ��
��ؽc,�����9�g�*��G�Kb|�����>�h����;��=��}��4]�9�ԧ>�s[պ`M`�_����ó�A�������	�yz���臞[a����RB�|<U�g�O��_5_*>��둋:�����sO�^��Գ���:��#���q��M1�F�i޼,���V��; ۴vj�9�O�z�X>������qg����~I_��P���u��t�g��.t�ƃU�S�ϼ?}�]I�M����N������Ƙo���ƴ{)o+;�ǥZ��owǣv����ǜ�2 ���9^[}-n_qD��n��L�5:�����l]���X̕�x�$�S�Ww�	t�ŠOt޹�W��9
��q������_���Z�xާ?�a���}�;�_ܑ�h���ŉ�q-�_+���p�}��a��@��!�ϼL��	?��g~�Gfj�2xX���Gv��n��6�9O=��I��H���N���z'���V_�㙽��e�O��:������x�=�G����@�+�UqJ�Ӟ�W��5ߋ�و�ٯ��!<:+�� x������Գ�Kޛ�é����;��c)��n�����躞���dӬ�u��la���vNS�ϥ?�����<������-?W�i;bS��<R�e�⒢����� [>|@Q_�����1�������>����ݎ�j~��r?U����O�:�.�W��s'�ܭ���YK6�+{x'}$�2���}�r���x�KN\�1m���6oc���C��.��N�y�yW�G4}1�/<�5I�=�]Q����p���c��ã��!��3P��*�i��fq�{?���9��n�+xe��lʾL��f�<��>��b<����������8U�_·���Z�OU�C��|},���?�|ܫu_�~'|�\���E���l��,�D��Y}ǃuי��Y�OW�]_o\��w�W�9������+��6ݔ8||�����P����J�_��T�fx�W����`��yJ�?�����[�^�j�U�W�������z7Ę�_�?58�w,��Z��;��1�󉫲+\^��NO-Y|�����7<';�2��y�5?F5�2�'�����7*�8�����zX�>9`p�~������V��8��
����1�o�E��G�.zSy��,���,�?���8����W�����ƭ	x8_@�;	�y���|w>��eX������+��_i?��9��=|��hx��¸�$p�=�	��g��߈!>���Yl�St��&��~���8[=K�c�e��<9��s|=��ڙ�=9%^���$.���C�~E�w>�O�1?T󱺟����Q�{fR��7?~�8���o�|4����1>O�V�yi��P�*�N�Rm?���b��r�v��im�A�������M��~6�go,ߗ�����|"�����B9�گ����/���8��2��ّ�sz��2U�d�-��Y��iv�U��1�e5?R5AO�$���~y���o�g�kz�/�ڳ�{�:�n�����;b��:8�)mb�ϧ�{u�=b9�����ϓy��gQ�{|��	�˝����3���<�>�9��[l��>l�3<�O����O���{�*�?�';=t_���8����z~!Ӄ�]�簪����Rف����wb{�h}=���zB.�}��oѮ�8�A��,S�V���/����f����$�[c���Ok�y����_?2�?�t����0<U�����y�*�z끑��"�����G�ktX�=e��o&��q�.�/Q�O��>k}�6��+����A<���z��*=X�O�\��p�=B�<2�X|���Ջ��qvG��M1�Þs�?��I���~�/�2.�9t���E�~C,�s�f�|�r~���I��|�K�~W�W�`�������	�wf<
u���5������ʏ���s�Y�1�A���Y���_�>o�����?�9}��o�v�ĦS�k)���_����wJ�Ƴ�vx�$�/��t���*������;�Szr!?������q\���|���,�}m�^��T^�0bt d�fo^�X��քˤ>>�˷�8��ɫ����w��91�^u_��k�q��S���nB{T>w�7;#������6��N\��ڞW�@w��?Kfo�8?�����<���+����A�_�i��=����yx&�$�}�4_Y���פ~X�sb{��ޡ\R�~�S�ǅ��r��ڇr}]ٱ,��8|������|���f��{�bُ���v��?���}��m�=����t��w���vi�˽3N�����F>��������B���yA���b���nh~�}�q�z�1�'pG���N6����1�%�*���o���Uq>��r�%�8����S��a��?ߏ�q<ψ�y�rV��e'��¹������<�Z������ǁ�կ�L��|f��M�78�'n�3��=��	6�'�]�މ�k\�˓w�~g��*����zy���o�p�?�������vu�~��*�T�g3~�q�ӟ����ݰ���ّ˥������	ۺ�^U�ُ̋��}q�{yQJ{>؟�ct]V��<�{I󌱸\�y�}��k竊?�a'b�s'����O1��R�],�s��;�KT��g+����_�ܛ���Y5��z[�_�����Y�7����~�x�������X��g�����c�J�Tp��^�ס�i'��;����T�1寯k��n�����e����������{x��3�<�������o�����s#��w��xQ�z�m��	�%�M�?����g��̏���go���J��xѿ��"������Y|��u�>e�t8�+����U��꽿���"���ga=o�*=��w��Z����l����v?���@Ҟ������Ag�w��������EMŃ���bq�����]������ؙ��{}�gԮ�yB��� �#���yzi�&�81�C�������%���j�*=R�WaY����PS�i\�hO�*����Vތ1?�����U��������w�y1�w�K��y^��j>V��v���5o����&�w}e����<�w�}$��c��8��������C1ާ8Cꋾ^�?�ɓ�6Oה��!����r ��^�{1N��8r�h����k5^��R�_�|w��W'���l>V�;��U;+}�=z���-�z�1��z�GG����U��d���LٿV��s�k��u_[�U�s袣���	����~9W�=̅��g[��	ކ��|�:�����6;f�W�MZ�O���܇Y%�u���%����s"�~��U1�p��5���ג�g��/�p�Qt��xD����_+�`}���>�K����w)6{{6c�o������}@�g�~c��7�w��D<su��^������W,�����c,�YܞQ����'�������ot~�y9���<?�e�ҍ�Ί:�F����p����{�O.�ϗ�X��ҿ�lc�S����W���sc<�����\�_���s�Z���/���gt�8��c�qY��jP����G�ϋ\�y�6�/��7
�:������7�~�_��ߌ1+ڳ'�ϯ�j'�g߲qQ��;�+����Ə�Ϸ}��}ك�R����/��z��+�/ߧ������>�?��3���Ǔ�^=5ry�Ӻ^����Ză\"��iϸ7{]?���u��݈�9���Wۣx���k�v���_�ͫ��-��8�M��k��|����o+<���~n�d��1�P7�p��*=�R�B~����k��%x�&�'�|�1|qf���lh�3�xW���dq��1���#^�\�e�[��`�C_e�m9=�m#�c@���=�+��A|�?��>�C�޹1֧,���x�܃<�x��e����N�S�w�M.�����~�	x�����դ������|�N�kS�V�{�������韵O�_�}W�M�՚\���_��=y��,���k����7t�l]��X���z��z^�ts��s4�7qKX�C>?5���߻ٟ�c�ռ|j�^�v�;�?;G����(����w���w=�}�3N�e�e{	��|N���kOo�6�؆�9R��
��������������w�e�����k��;��?Oక�@l�-],�G�����	�v����}��?ݮ��U�Oو�#�m���N�����b{ެ�kO�x�������}$��5�O�d��{�8Ng�Xγ8?������ɏt����q�9��\�onO���5��\{/����e����#e�{�J�*_�C�_e�O��Y��O�1?�\U{�e��pk��G�M곏��M1��׿a�3{F����a�2:�tkޑ����)މ�&�ß�E���~<��r�hO%7��L�(�Sz���,nj�}��'�'��7���aV���x*̝�p��Ƥ_�Wo���,������\�?�������(��9,�b<���A{�^�V9�}L�/��V�u�A_k�־t��V���߮���6N�����]��I}�WA+�{?�'�7���O�tc;�o���Zϩ�����"�*l��"�צ��~�J��$+9/��T���/��3��S�󜧏����d�S�%��g�Wy�}6}:{���9�����>�gw���E��:���^������>�9:������ï6��>�+���ܟ��<~l��#��;�,����Y߯�����9��^?���Y�m�<B�CI}�'�:N��x~�WX%n�!l�I�����kqF~&�7��O��������?�D��>%�g/�q�a-����ޟ�����UvK%�'X3d뵙�u_�I?C����T��nG��u?����/��cؗ��U� �ϋ}~����sO��}a����ۓ���-�P��x���v�|W�'b;��X�����v����5݇R�@�=�}�w�e�����;�z\qdp�s:�w������)p�� ��4ndC��{!`�@������/g�]�=�?���,yoX}����^���"���yg!�2{�����3�������c��P�C�s<�~>�7�#^�?Ttֺ�E��6��Fn������b��8��*�V����ԧ��	��{�/�q_Jԁ����������wU�����޽:���q��3b�?_�?���	�L/����a�+>����[�|�����9C������Y��~��E%?u��~,��0�`�~�Y�(pʓ�\6�`>#���
�<��U�|�[1��-I�l߇4��a}����_����˷�^�|������ϻ���4ToM��>,�{����~���۩�۔���|��c��P�7o?Q���;�G�w��]1���n��=Ü�o�v��kVm�^o��g?w����[�/�/�Ƽ�?����b�T����{}̧j_�����bD�ٟ�fÏ��<��[�_�+�����v��}W�O�Q�7���N�˱q;g�@�g$x�>ߊ���˄��\oc3��@|_��
O�1�a�!6t�"����s���xĲ��Nīh~-�oW���_�e�������y�b� O2?��s7�|U��o�,�1�7�����_���O�ӈ��]�_i��w<<���(~?�����&��։�~�i2��_|k�����h\�չ$o��]�[��q��vj���*���G�;�*��u7��z��U����������L��q��V�?�گy��#������Y�fh��Kb��������	�y(�ә߹���1����a������W�U{��f�w��ㅱҸP���j����c�wgi{_Z��r>G<��X���C5��'_^c��~����o�s4�n�������	}6�>�������v!l����o·�Ϯ縳y�Q�a����M���aNb\>����kY�A��~�Kޣx�#����ݞ���嵍Z���������;�c��i����q�7��q.J�$@>`�it@~6� ?�uA��!�x`���X�gJ��I}�g���WS�X��N~�)�����uWr�ãtPz���s��?�~ �O�c(g�?���0C��#1��Oo�׎��]l�<ϡT��p��;�x~}�ÿ3��S*���t�z����g:<[V~�0�f����[ٓ|�������ٍ_/�?�i���1;����l���j���,߉��Y<������<s9����YМ�����'����)�|�{s>�l߁� �����ߍ6"��y��_�뿱��
�sSk�G
��N����1�+~N��vc��z�����O~���o�{u{��[oI��r������!.�۬��X�[*9��h���̑�9-���怎ށy��]�G���ٞ}c<��Dn���7�����noW|˲Sܸ��.�s�椾�c�a`ӿ'���;��|�������w��\r:�m�{s���^��~�=�ῡׇ�Q�R_��vs������=s��o3�!�s�W�0�/s���Gć��tޑ>���/i���������Kz=�zz>��ٲ�'���\�i�n����/��h��=*�]w��Wj��}���>��b�o��;��&�/���i'�_�z�ʆ��_��u���.a�'�y/�̡xM�G�K�Nq�Ο(>�#�K�����}�9O��f}�����g��� ���u�^�<9��*��[���9H���t�S�������9����ĕ��28��V�_�����;2�˙�_�]O^��p~���Nv/�g�;���p���K~C�NL�w,{N���'���(�{+��ƾ&�ޟ�ߍ��w�W�T���/]�IEϊO�>��M����K;}*}*?C�K�k�g$��?~߄�������y�����<�vu�0r?��wk���qYgG~����d��c���ƅ�����!�TT��ϙէ^��ڳ�5������������|]��}���y:��4����a��������:�|<����sZ�����ʎ��1ֿ��{+{�N�}v\�B��G��=4��g�{E�O8��H�,�W��]����9�<�������|_�=����/�(b���l�]��]��������z������w���3<�G�旎��D>kQ:T�F-S�~����v	<��@�ȟY������D���B�d��<?��y����+H~������We�h�����ځ�x����}Y��*;jU���G�!%l�oN�Wx���kc.C�{��j�7B��|S� |w7��G�uqq�|�����}���^��f~Eꖩz������'��=L�����8�+��q_O]ӟ��&����J����g��o��!|@�)�%��ưw�T�Qٟ-kO��U���j�G��X䍟�����p��bW�m���ע�w���ߒ�b�sv����]{�S��݇�z~���$�&p�	~���؋�Eऩ�߆?
��{��u���~C���8�	��{���~�wnk�E �E�n����B7�&U���|�}���a��*�B�:��a�U���%_�w�����:��>�W�`��z���%����ت��-�u�>����]��X}���n?���,������e��
��u�*t?���9��_����u�)��f������������T��q���8|�sV�k���C�G�?:��~������\���w<gM��;u]��Z_�K+_U��u�����{���|�y�>�_��1�g�ᛑ籯�s��;�i�x9~���4��NV?��Z�����o���5�<.����B�o�pF��6|��ٯ����ԇ�torc��+�:�i�>�N�����9�s���g�-��^��5�W�O�w�\���^�q}�vvy������O����p(F�{���t����;0�Y|�ׯ�T�dq��~ �t;d_��{�z��3����8��h�O�`w�.�7�"�<��F��J}�sc~���<���~q��{��_��c��Ё����n~��[f���i?�#�z}�����bLO�Qy~Ut���W&��~�>����{zu�]Y<�<�}_�k+{F�{;���L��c?�o��mOf�����{{�܆�a���A�}��G����;~���d�)*��_�{�>c�֋b�V�ٮ��~���v8��ۓ�\\����|��#_a~bU~Ҟ���ZO�8>������	~_?�}�?X�|J��,���I��O���Z����������KyC,�x�����cp���� x����\���r �䃝>Y��~�)p}/���W���|Q~`�^�?ksv$�u�G�>�	�|.p��\�0������?��^����'r����Ng�_����< p��~~pKڟ�_��;�`�{ܾ����XN�.���=�߭�ζ�辆ֿ�?{|��V�OǶ��{5^7��C=o��w:T��5���ӟ��~�h�3�������1^_Tq�պ��E>�+�_���4���7���ݫ^����;��.H�n���l���:����aGb��ʈ��UV���x������<ƳO�Oշ��0��e�'�g���c��!�|��BN;ߟzj׻G���	�p{,�b�߉�5;�u��ݿG��|}�<��/�!��)��e:W�C�O��g<���g������7��������p���1� Uy�����`��΀N�s.�'�����l18�/�������:�f�̚^X{G���}�=����Z/x��ӓ� ���G��u��mca�����Z��������W=�����L.�^Ӓ��|�i]���d^�K��)��F��Bf����}������y��?`x�~��ύ���g�sg�n��z_���Wz�váqg܇{c,��@�o����^P8K�OM�O�ՊO���ZrrO������ �����g�P�~]�)�����b�@��M�O����wCV8��1/��ϭT�e�׃#�c}\��K1�$�W�z=�U�¯�S��_�k>�ꞩ����+�|e�ͶF�ퟀ�8�v�*_�Ӈ�9}�\�[��y¼�C��׮0<�k���:�qߨ���v5όe�~<���U?���p�����p�0�j_(��/�y3������P?��#���#�>��m｠�z�|����6M���߁N\N�J����<��j����G��y��>�����*�3�~���������Ƿ\�q���un~~�����l^�_���ɫ��s��`/�`,��;:1����w�~|d���I�����{;�?%����H�/�䞿W������>
^o��+b�O��E�_�O?�k��l�$���*�/�Ը�)~��.r���ωAn�}�{�l?�9����q'�G6��������hC�ɷ�ޫ��8��8^��7�LN���S����U|q�_�s��OZ�?��?;��ɫz3���}��'���Ry�p���G��SC�@~g��,����'[���q����0=�R�� p���l?<rQ�N��u8�F�t0v�s��1�>�c;g���w����
�/��J��|�h�@*�Y|�Vq5�W�Sޞkp�[f�F,�g�O�:W�k�I���x�?(߲��OO8��X��_��a*:��&rb-r�|,����Ig�W(m�~������>)x���*�[�f���9����஽�j��5�i�;��&����6����v������?������4<8o�G1��K��F��QK6�,.�|�˲�]�p���v:�y�W�zX�)��֚���4����zM���GϽ꾘�[�u�Ӈ��(k�o�滞�9 �����j7��6�3���鱸�p�����yy,��!����7P�[�����<�gR�!�Tvr���5�w��4�L�YU�p�����Y,���Ӣ�T�_՟o����Vc6��}����֭�����e�k']oV���������W��]��k��i诚�N�j�=V�u�gEm�f����|
���s�xҞ��l�Y�ŧ�����N�zi^}�3S�=�r��r1��Y��q�Ʊ���_���	���A����Cց��Y_����U�_ٷ�^��۩ֳ��m����HBεUz���K�����b,���?��a�m7�Z���րG�=4�"k��UІ�Ý�����0�$���������}��߀�q��p~�~�]��s��3�[b��س�͂v�<�o!�qFT�i�?�_�*��W�+���,�o���ت|���ix��?{^_�W�|�������~D-�o�/�.��],����������<X�`��1�kQ��d�y�l�V��=S�s�y��?E<�(��T<�kM�V�k�|bgƶ[�Ϲ��o�w�7��V�-O���}U���1�O�>U��~�l���ec=N<>﴾����J����q��E�7.�|������u�8��En̰^B���_���{�scl��@�{$��/�_��V9F:������z�a��w��5]�8G��o�;b��o�e~v�3��X����{s��s��#ͬ����u���+=���/�kT�؍l��_��r9���������=M^�^��tP�7h+��t�������.o���y����z��it�]�B�'ʇU^V��k����/�slo���8��{A���e���F���K;�w�8~��J.���:�}B�%No��@���D�o~N���^��oFΟ�C��W�6�����8+������9�wy�R�w�M����y���i1m� ���O�o�!��
�������q��"p�Q��*���tV�A��zS��)��.��N��v5搞g�i�q'����u�Dy�vȱ�n���~�S���d޽.�<$������ߟԯ��/�_S8��Gͷ0�n��Gb�w�^�|t\ˠ=W$�3~ \�{�Skg��?c_�{�\R}G�����~�.����1��he���,;������z?t?��ϯ�����_}�s��Ϥ��1�9�}�[HO|f�d��a�m�*��M���7��Uȇ�1�s�T٣p��{A�:R�plWэ�i|>���.E��+<�|��#�m�A�Y\��v��*y��O��oο|U�����[��oj?ic���>?+x��qe��1��}a����0.�'��{�տ�ͯ
n��޽з�|*g��8~?�瘴�������]^��bqW�bH��S�a�}��u�*}Z���y��W�]x��v? ��gޟ�n��|�V�wޣ�v�%1�����s �_"�Ը�Ww��2go����j+�<˓����U�Y����=�툍�毯��t����b������O�oYC����j����!��C�<��\��<G��f�Y�΂�f��*��7�C�c�b]��V���!JO޳ ���&�O�����f�"�q�j��R_ۣ~Q�?C��oi�m������;�;k��W9�����������5�nx���?u���=;����D?T.��i�^����9t>�|+����E{	tV}��^z�q�����t�X�7�\@fW���C_]��w�ռ�Y�ة���I���q�|OA�}U[1�:h���@k�gG|)t	���1��n8����R9\�*��)���/1n�Ř��U���Z�y��Ը�����3���=�{W�Z;�8��nE�/6վ��H&O��J���Y��ޯU��|����U�N�P��_���E����T�Z�~�� ���Ʋ�>R�gĸ�¯��
�ҳ��E>�N=?N{7�c��4J�ʯ�y���n���`C}y�k��P�����ym�?�� ���S�:^U��N�ɮȟ?���yE�ݹ/���^�9�?�� _��K��N}��v�{n�����C�-[������vx����#Tgy <n��+ۿ{w����{��;��+p��8.�)��.�h0�Y�+��N;�g?wI_%ڙ��N�����gu�)|��uo������؝3������|��Y6~Y~~���`3����X�F^���P�Ê>u�Q��ps�Z�k�C��1�o�����K�#��s�{��C~�g�f~uC�#M�^R������8|�ൟ��n�Ut^�w��_9?�އbX�较❲��Y�w�O�YN��;K���.����U�1v�3�����v�N��㸸_�Z�Q�y�L��.���a��w�o�B��pnE��7�S�
ï�yJ��j�����Ǹh~E��+�n,���Z��Y{�N�*���<���ٖo�E|�L�69^[�΄.Cd�	��~�1����r2�A��j��>��~i���-��y��@�G�KV_ǒ�o���_c=��~���y���Ÿ�n.g��L��|Y��s��	~��<��|��D�7��Ul����7����v[�Q>��P:l�� �u�b]��=d�:������w���[�����|�>��o1J����L�7�|t���o'b�W3��bp�A�[��N�C�{�K��y��qV9sf�y��=���S���{Y��N�(�g�>��j?�~[�3��������8����;�[e��=�͆_o�q����3V�_ı�S��_����/bq?�V���o������P����]�W%��//4<��G�[�n�����]��yG�}�˕=�8?�B?������ʟP��h?]f�ݔ~y�I�[���?�硢��b�xpo֔�{��I�Z��.��_��(�T|�z����Řo�n�_]��W��d1�;��E�sG��Œ�
Pl�t��X�gY��yq�~K�߹����&o�1�h���a�pܴG��E��߈\N�|>�����<���u.��1��8Nf�c�qD,���p�wW��7+�.�oPg���N�C����sQ�w�,N�O�� �S�#��#/�rNݶ_���c����rw�R���͗�����j�����WJ}����o�[�o��Wg#�������c���u]�wθ��;�P���׹U~��.?�ƸN��z�y���vle_��3�L��x��\?��yW%�M^������ig@)=�u�+aޚ����h���������*�djހz�ό1�*y��a�/���pį,���h�S>����n�v^��?(0m�z]e�����%�8�J����<�x*����;:e�ݐY�>����_���,_��o"��o���ZL;�O����֡�_�}�F�7�|�a�鮵��e�������7Ų����46"燝�se��P,��>{�M�3��J�;��뼮���o�Q�{�+��ʟO��a�t]�R�7�|���C)='��}]o7�@��sy?#�cU�I��7��C�Y�JT��ǝ�|�Z��e��a?���K���q�=�vV~<+��cȋ������󉯋Aa��Q	�=[����9��_�m.�tP9p�������c��EC�٧	��rj>@��w��_.�9O��I�kry��?c�k�}R��v���p�@,�W��,�9�`��:�3{�+b����]G�f���w��z��s<��y�yTX\ϲ����y�S������I����Ox�������ώe>�9��/�F��}.���?7r����Y@�[�k�'�u����#8�v���~Uq5����s���O��.�����f��������C�fύe:{�Wſy����.Wu����;U|��Ot,�ܗ�忪�����ۢ�W�cJ���U9�ͣ�b̟������f�S��5n������j?�e�8I�W�(���}Ʃ��(곞��q�E�/����(���:}K����a��J������y��^�O���b�/��0]WN�'����5V�ߋ5F&����5����;5L�����{�6��|;b�������-KƇ�q���n�7<�y'�,i������s��'��������s|n��I��o�_�y��T����}���L��}(�����U�/��<_+�J��{uA���9�W�x�X�=����n:�2�����\�k<��x�^����°'�}(��{��?���X,ӭ�3�sXc��@���uc�h���r��<��J^V���l�����#���X�����sİ�0�7��_���B>�~�.p�.�c�Y���{�ѮW	��c�o�?1�B���/��W�g��<ي��۳q��r�:o�v�E�|�i!kϚ�֧,�g�
��⤾�뼦�/l}���)�v��u��bXGj�9�\�%�����������}m}��\�#�W�~����=�s�M��Ƶ����K0w�۷�O}Q����d�;�-G�34�������Y��k��6V3��<?��yc�r����
1,���������j��ʷ@yt��U{X*���߷Bfi����)_�#��~���w����d�=>V�w��
9����?b��Y}�C;��_	��|����yT�GC^�A���t��Z�~��1��l�P�c��?�v���8T�[�,q�N[��wa�<��7�d�_�?�����(��W���z,�7Vy��U��v����k.��s���l�9k�v�����������\�G�9������*�+�T���V׭�����P�oa��#I;��h����qW�ۺ/	�؛��_���C�ն��N�k�j�]�����7��{��=�X���O�5�Cv���ƕAFj<ؼ��opyl�YZe��>/����8}V�+��9�9�q;�on���w�wM�/���/'�E�6���bzɾ��*z_���Ov|�V�+�vfo삮i�ٻڟ�W��5�5�s����P�QY������R�����9�W�g���9��mF�]��r����}:��<o�f'o���rx�E}~����q@�e牦�{Y\����/�ݟ@Y+�Y�UXs�������V�e�?�Nʯ�Z��*�����|��ħ�`c��>�>������4�~]���/r���]U�d�T|[�U���^Q�����`k_-p觭�Cv��:��t�MqIwu�x�I1�+�士�*?3䶎#���u�����������>S��U{H_?�3}��a���cLg�W=uo��p��t�m� �ω��ߛ���ɵ~&�g1��+�C\�c�o���+��6՟��?۱P�xe��{�&�j>���xx׻cq���O���8+Ҭ�2pǳ��pyB;mWL�7 �>��>�cp����	�g���A�&�u�����2*�7aY�W�9 �a߿^�we?Gr$�{\ݎ�*���V�J�}3���}��N�~����j��G��l���v����/�95�7s�:}�_�n������c�A?�4�ˆ�y�I�w'�!�w��¯��]��x@G����Mh'�s���΢gg������_i�_c�G,�o/��܊����[{[5n��;�]���畽��\���C`���gq?������q��/��~�?��v��s�����;|5�L�g��®���.����P��*�z�����X��o�c8C�!;�l��/��9���ߕ��7��
�}g� ��/!��<c�Z���7U\�Լ�����@����*j}���sq����_C\뭱�'1<l�z��Ai����t�E���������Qﷺs�c�����ځ��hc�9�s�����?�\D߭��~8�;�� �7c{�����U��utiq;�A�N�T|���3;-��}7�	=������>rc�r���*}��X	w�ڸ.b{��ԑX�������=���g�x�j�������n��Gb�8���^�����'�?�����b�^��@)�a�$�1;����<?1���>��
�:b=F�zqF {P��m1�?~���#���Uz�|���ώ<��3��Z_g�1����T?K5O�n������?eB;�(=�N�|������k�/�e>4���<BM�~1��=���Y���L�#}�ғ>�_��_��Q�w*�}�8��t������?��e��5oX����q����+����	�xE�J3��}c,�=����s�فb$���GT���
�s�
�}�ل�MG�~�}����5yoX}��~`�|wU���C��c���������׿!���wʷ������o鸿<����b\�󕏱�w_Ǘ�?��K�1�,���}�N�e�?;�����l�����8��#���5�8�=��
���8����W�8����T��x�����f!W�Yߛ͋0�����N��}�Ӓ�����HoS��U97�|}.����_㥵�:��|�EN�*og�/������<�����|5�w�:�>�-�͞���ua���m����_T��ڧ;Y�'y���j\؎��}��,�^�K��Ϟǉ��K}���ok���ڪ+���?1V�����O���Xi���������OZ)>�Hڟ�$��c����g���|\`��?��]��0<��T���<�������1���N�,_AD�s^��4?֪�]A.���P��J���xA�G�SS����~{h�c�A���Ɵ3�G���h{�9���y�����W>Ay��m�u=5e������yw]�wV���Ά�h2��o�3��Z������Sb;�X뿠�C���I�Pɟ��[�|7������`]�Wx�~���ik��_Ơ7������?c�{+x����]�K{�~���݋�3xE�3��Z�qJ~ު�W��b1�z�e����u�)��1F���\n�ڧ�.��)�~���)?1��pټ����=�q�%r�������X�I����<+����%�΋i��*���E�����Τ�)���/i��>����0�6�����_,�ν��X}��>��˃55�z���{�w0�ͯ��g��,�~O�k�3�W�3K���w���Ƿ���K��j� ��{��_ʹ��N����}bl��7�kM��=���/c<^��ڍ�C��b�z��
_�����kU!;�7��D���T{���b�$���|[�I4��v�T��z�ק�ۊ�9G��7��X1�����b��m<c������#dl�,���w�[��������>!��'�;�_/2�ԥ�$�ǘ�x�v��9��u\_$p�w䫳ϛc�~O8�Qv~�}��q���<:&p�۫&��|<Y�,n��C�mn�7�}�T��Q;g��Y�e�2���sV��e���8�h��g�x`mgu�$
�)������/���:��N9r�<c��`h���uyk���e0��X���7 �\_�tНw�g���k�O��3c���ϣ�d<��G}�������,�����1�W��G��c<��v�׷&~V�f:�E��h�^�2�Z�v�����=*�#�O���/�W������Z��S�#d7���E}m'��b�4_�ѡ��Y���z�#1�>�i?���o����|�X؟3]�s��F�g�i��@�_��c���/ʟ-�/�����o?�]S�����S�0�G:�7G{E�����M����&�J>�N�j����%�����_�F�ίy�_o��W�_��%r=�txY�'�M1�2�|��g��=��3��T:�?�չ	�7��Ü����ON����ޏ���n��:����Y,�A����2�]�_e'?����=��c���7>���u�6|����T^�h�/�y�����y(��OnUa�An�������W�-qj���ǉX��+�;`��T�����]?j�m�ϗvb=��k,���'a�����v� ��k���<~�~�a�@�
:�>��x}��,�]��<�;���
���e�\/�����������gc�(��U�?/F��t�`v���1o�a^��w&��|S�ӝc����X.q=���U�焴/��c?	�	G�~e׽*�=Q���y"ҳʓ�r�Xl���>��;�v/��q��d�sʅ��}i{��ۃ�a�o_ֿ߾A�����O�p'��R�OJ����O�Ϡم�=gx2:T����:s]��gĐ��S�޹�K��O}T�y�(��Clُ��~
�9����|����=�y��ht2|��+�1�Z¿�t V�U<�lL�%M8�Y�3=��{�ڻc����q�����v{��v8��>������u�������Q���w<*�!/��.�}�������5X~̧y�~�_�MQ ?�}՝�ᙜ�w�?��.�����֞�������u^�!�㡟nj���wܯ������(���9�����(�+��]���H�������f�u��2��������Y��Ƣ��>��5�I}�{��Ϸ�cmڿ9F�_�(պ,N}��,�?�8|~�v$ָ~����s��=���{;�}��|^T��*^t�s:�7�7� �7�=�����;��=Kڣ|���V��G}����á�����B���W�˺*�u��~7��Kc��|\*yE\ʇ,ʇW?oR�G���ʙ=꫽���������?g����{���cOgk�KӸ��?Oy�K�[���kT�O9�y�|���>��Wx�wX;�v�>|5��J�=h�zS�aT:���c�L����Y̎�ᝐ��ۺާ=��ǫu\������־%r>q<�
��7k��"�/p8�c����d���7����������o<C?�X���q:�?��s"��W����ee�wʛ4�a9=��I8/Ύ���K���}��<���Y�g�S>a?o���dr��깼��Mom`�����;�����
���?��b�U�<�.����7c_ݟ�tP:�o������uS�����\ѧ�����JO�{��������y�OQ�:'�����Un�|v���:�Du��/�bg_�T�R� �M�eWzY�W��^�)xN�O;կU�Govח�߳U;��9	�JNz�����>y��'
��,����U���F߻j��p�،��E�0�a[�z�\W���y����G8k���`�`L�;zN��Wz��'f�"?��3؉�����v�k�e~v��X�b�kB}f�����\��wo�ʿ1��{[�LTr��ݨL�qJ�~���|���|�����h���%�O����Ƒ�����������]{�yJ;�ށ��n��1�'�!�����7v��������cs��S׹�?���N�{]P�������1�C��V��_�=P�����ř1ޯ�\F>1�OO�pn^�!��xQ�S�<��e��kS���U�݈�_�:���� �8}��N���aa��+�V��<Ng�9��78K������-1�1h�6�_����?�>��.��P��[��3���z��Ϗ�<��.H��*�����h�0V��4_K�_I���a�f���d��T�
~@����+{��_�����X���9�y>?0��Z����Ժ�o���D�o���9��q{l���������'�-p�+�x�����W�g29\�W�>�'ao�����mM�������~,�=������c	����8��{D��I%7��:�5.Q��7����k��c���5?C6��%tX�����?.�����?i]�N�����ƞl��C<,��N�sg,.� ����gk��-�:���9�J���g�N���G���g�q�x�,���;׉~>��y������8�#i���_]��5�Yܹ�/��ݭ��(�1��[1�u��+����|M,;�g����3�t�<�c��h��#�G&.ҭ���ك�[��W�=�~���o����Z�q�h{��z�1�?S{<�W�2�Eh�����q�g����\����,��g�uċ�7�"Vi帳��f��`��i������|�����	���x��iTv��u!K����;&p�q�=$���LU�mO��}p_杞�C9;�C�����"[_���������>��a�3�~e'�8C��C{�\��bD��l_#[3�9����I���q����q�zN-��Gۯ�/`����Ύ�u�ʇJ�h��)ǜn�>�֍X���g�u��L��W�N�<����/��_j�>
c�	��zP�W�r�!�x	�oD,˥��|�~�Uv���B�|8>�xQ�ǥWy{���o��?�3S�
�3��\��~�v�^��7��������R��>����{�����>����Q�O���J~R��>S�*�g����zu�N��cXw�^����+�V���x��c~��~�_�i�S�7����}�- �w��\�=�]ϼ�ul�ko�܏�7���b;<�.�����A�{�T���k|>�C{�p�?A���~F�9d�c<{x~��6��qm�����ó�h����&W�T�Ӕ8�U�w��t�O�sƇ�o���8�>=,p��`�]T��⓽���A��|����k�=����uÃr����V���ໃ�?b�����l�g �1�:��j�[���o�q�d�{��`���y���E���߫~u����u?;���m�7�o�e'�kF��П�t�Y�>Es<N�1�}����޹��\G��9�/r����k���y��1ůr�������!.粿;i�<�z��Ϣ|v'x���j]�:��2�����zU��N�(����k=��b�U�֧|���s����s��io�����ĜV���W��|MG��zR���[��w�#]_��<���z�e�3����~T���8�h]L�O�~�ۥ8?1�T��p����;��x �s�> �d�Ur����ۿ�?C��2��7��T/��|�8[][��Ւ����p�^�+W�+��T<Uܚ��>ER?����C�?��C��������.�>l�	����G��;�A[�3�s�Y;Y�s7N�U|^�w<�ְr,���	�n�%��]��+��gv��KQyB}����i�����T/T�Ah�j߁��`�d��j�fW��5�ׯ��Wz�	���6��]��@K��ۇ:~������@�k�+�����x�Sbl�О�<���},ν,b�B�Kv�s���9,>.�{\��Ł�����։��`,��_�#�P�O]�r	:�Ԥ_o��w�FL?ϥ|�z���}�N�������\O�7������K����b��4?y�����Ha�d둝�](�i��8�m^�ww��jx����9S����7������,o����vc���k���B~���1ȁ�NX�����kX�ܖ��Ǘr|#j��α�~Uz%;���Y5�=�1�,��}u]�Ϊ=�^�X��g�x^h����������\XG '�7Mh�v�x��ϓ���c�#�oO�������x�gNi��x��w$���g����]�L�C����/��_���z��Y<乆gO�s�?���v��5��}�ʐ��y�Sc���~��bY/G,���\�s�]֯�O�߽����-��ߨ����q�^����ox6����=�dyw7�n�h�'����w+��t�l��-pI,���'�0�~'Vq���CI}�U�W�qe�Q�U��%=��C��?�?�������^��S��K�O�g�ϵ/��N&�|�����C�_�������i3�G�?�3���1�I"\�S�d\ڨ�Z2��<�w؁X����V��6����y���s��{�����;ߏ������y��~������/8ߩ�v�O�E�����L���]�w���;��:��}�O/�L2�M����l��?�aofq���*N��0��1-o嶏{�?Q?��ҟ�%�k�?ٹ]�����#��1���z�/��A�������&闷G���ҡ���R��8�[;5��[ǔ8@m���}�?�~m{�4P���g���(ک���q�R׃䫩�]�Ӱv|��J����ժ����/�1?CO�gp8��n��
k�/o���ϧ��N_�1ֺ�Y�P'��}K�O} ����
*��}�ST�
�u���:�n4��x<O5����i��w�sI���������s��u�2<�Gq���?���U��r�tw���v�T{�i��sb_������m6�Z��]�xt���y���n�/���1ޗ�����s��,�~*�[�����<�� ����X�g�+��J�r��1�',.�o��B����������w�pQ�'������ۧu�۟����|@��/x[3��ψ�z�����u�����������T�'_gAf�7�x��a[}�rV�~S>|pl�@Q�������ոT���� ��w4� �{�Mu?�t�M֞�N��ݾ~�x'oO����*����Y|��y՞j_��e�������|Y��=��Pcp��91��|/ک��aG�8��S����ڿ8���>Ւ�i��κ������Q�$�������X�g�U�(����A?���)m���>�	��:M	�~+�+˯�v·bXw_ߚ������gŘ?)��D��8�q������a�/S��y���1�ϑ�������iE{�}�j����v)κ}vQ?[_�=Ʋ���k֯��ߟ��x��p��:՛���o���o#��s��9�m��{����C��@��������^>�����X����5�W׏'����Ϙ��'�<ߊ�ȶ=���������E�w{�����ߡ�$O*����F�+pЋ��<��{�����ď�5.N�M�W����[*����-�ۦ�fXo�:�W��}]�p��<z������~ʔ���vؗ�����}1���Y���`�h~��>U{Έ�;{/�P?�;�[X}��#v��+�#����S������8/����9w+�dq�N7�S���@(�V��1��ƈOfȽ ���V�+&��ZP�m��$7X<^EK�_�[}�J�W�������=�u��G�ׇ_P�G6�.[�N����ڱ�;]<o̱��z0���Þ^�������XW��N��b�ǘL񗲸��T��Q���c+y�����S��'Y}-�;��6����w��[ ��霂���0�j��}�~�g�+�A=��M��'b�zB�����#Ke�W�T�7[�(�\�H����x�D.?+���ͼ=U<I����b�	z������y;������<j��7Đs{V���5���⾀5���핟�!w����T�vp]��8|T~�}~�^���?�pu��s�/����]1�!x�U�<�7�>�T~ޯ5	�ɰ����y^,�{|���Tk�w8�ަ�鯾K�ǝ�����݌>�{��sغ�۰��>���G�b;��*��w.g*9����Ve�O�!��#c�KK&?���������rށx̟?{����������'��}�yl��U��'�� �n��G�^��������a?�_���,�_�|�Z&�.ڮ94���by�#j�^�sO6��4w��eոWp�E�r�]����3���C�y�kh��Ȥ�޸=?�[mR}/�]|4�v&���<�!���٣rO˔q��֧�닫<�ۻ<�����r޽8j>��<;�WV��Bګ���ޠ<=c~�������E�_��C���a�w�h|qVf�5�8粦qn�т��:���}���y������H�
�!U���>�\�0u�U������ƶ|ZE�����k�6�kol`�?��׃?Sכ�k��	9��!V�g?]�U熴L�oӎ��+�=�������^��>��1����{뷷�4:m<G�CN��w]wl��o��_��g꺯����c�u?-pʫJ�{O�g����H���{�/�e��~�z�^>�c��?�N|I2��39�G���T���T낯��D{_&p�5 ���;������by���Q�3�A�Y����R����?�P�:�:o�}P�_�O�|Ѱ�t_�s���x�=�g��bLg�u��g��H����
��Weϳ�{�����]��3�ѿS����y�y�;��M������8��xS����ϸ��W:(���]�)p�s���%x��\��8�>����G�|��^�y�(��������~�o��^�o�>������3�y�}�`C�K1�?]��_b�2��=X�#�`������9��_��7�[�$�X�U��x�Ѽ��Ҧ��Oi��=�5��t��X������X��Z�|�>pyB�P�)�]��G����c8��}c��E^�;t������>�-�<�I�l}�*����5[wO�)fM������� GfW������Gz;o6���ૃorvc��3�����������ձ�Ӹ�z����s�{}^���녳cۿ��R���n�����K�~�o~����Ԧ{��q�wy����Wzj�q9{ .x�gaGB�#�:��V��c�(��_.�ˎ�X/S_��:��3������S\K����d�:l���=�%=���|���Ӿ��y:�j~g�KY�Ư�1:�t�#��H>�<�{b;f��M�珱�<?l������篵�f�2}D~T<��Q��O_��>��8�G��XUyDw?��1ܕ�x�}���IY}ۗY�cE�����̯x�����p��Ze�w�lwQ_�|c�W�+��P���������b���F�Y�/f�!��'N��<����2�Sa^d~�Ŀt^�k��S�U���ñ�и}�Ƙn�������r�|�T�f���}��nq?5杮�N����*���7��~��>%�t��~�,�EuNp���ܟ��8~Lωk{����\����a��ߘ����#ꧩqS����sE\:������D�7�u}&�?��wk{2>-7��;�oO[��z],|T�7$���O�<���H���|p{��������$��_�{��0�r�e��K������Ύ����g����	�Bn=%���!��G�OƏ_��L���t��0O��5{��5�,^��Dn�T�Ov��Z��;�o�>�6*�G�*� g�{�wj���σ�T�8够-�ޑܫ��w8��,�����]���v���)�䊟YܯB:0.���Xn�|"�㑤�ņ_�8���y���D{���������'bY�Џ��L��1���'�׃���'�0������}�qY��S"���;����z� ��������F獿��Ok���c�y@��q��Q��X���Vy!S/�e~s�Y����:^s��ه��ud�|j<����8@�Yh��\�c���~�~�zy�}��=[��y���W���蜤�����ܐ��G:�?D���m��������1D� ϴ_]�W<պF�@f~��~���5�?��᡿k��>��:��}u��y�=÷�2���$���[_oҟ�g=�3Pͣ�����;f��s����|g��L]7U�W������S��1����:^����O�2�x|��z\��ԟ�/���<S�H,�����yF��c9���9�٣'�w�?W��{X{�G`^���.���E[�^� r�\�=�*7��s�.Ό�<�9և�x���xF�Ǒt9+�qt9��T���'������{XS�:�}�,��<�r%�i��69�ԟj�s�9��w�y?3ƅz�����>��t����#J&'��^�S��\ނ�q�A�C�o�����G�o1��n�Ş����wl�q�`�����Of��Q;�ϹG����8>��b�9�~3�m��b����Eu^��)���b/q��c�����^�qr&;o�r^�j{��Y�J�����7c��2Wۉ��y��q�3���1~�q�X�ߞ|0��F�;Ź)���8ޱo�x2��x��&�����tC�Q?�zl履�����+��i1�}R?�c.П�'k�U�g�ٙ�F���u��1������U�1�S�o��nxX���$qu��&{֛��}i{T��H6����T�)�)_\� 6ǉ�k�~|��X{������w�8����?�Ź��f��{�������������W��K{��_1�?���O!�x���`��}/���b�z�������̃�φ�v-��~!�m�w�}��x�ّ��t��x�\?�Էy�����]��~�yw�����X׼7�C�����E��U��)�/���>~s�.�����N�j+<�=�?ryU�M��U�&_6���΢�{<��Yx�]9}�>�m��s���� d�w-�׹���s6��o��R<�_ex�G�I{���Tv������ߴ����������W���iW���݆��>����z[o���~����k��b{>�p��x����ߩ� �V뎊>(�'��h���OX����q>4�w��qW���������K�3bo���k�>�,D���ץ>�~�v.������⎴~5�~�	L�I��}�*���Xaw�|ƞ ��7	��u1�˷\�)}~��>�,~uo�Ӎ|p��~�zz+��`��������"�S���a��#8�}F�Ǒ�S�/|��F���F�w^�a��@>�;��m�ډ����쪆��&��}��x���:�{:|��AqW���G�o�fo��c����d�-�����?UN�g�
0���f"�t��gӧ�.��ύ�~k�W&�2<��{^���k����̯�g�玸O�k_e�<�Ӏ9g	��tY��7�Dg�n�<_4ǟ�i�]o���v�8�?����8�`n������T~�l]�B8�s�~�q��yU�y-0�ٹ6�~�^����/Y�א��Q�)��M������
��Kz]�O�:Vv2�@��}�ΧغcT�����Y�Q�|w;c��	�#<7�_������-���R�)����k.��5��'���t�������#r<찭�)����6/�ߛ���OΙ^�����+����Gh~!�!��Z���xf�s���q*=��[����N������tګN����2�����c�^��)�G��>��eviE�����<}���L�[U������9P���J~�<S�~MG/�B~���\�λ*��Xה~�u�}Ni�86���=?R�2�s�=��U|ڽ:�F���^����}����C�Μ����{;y��K�T��ո�*�{��sۓԯ���{5��� �������@��*u���K�������'��z��;ܧ ?�N�����/L��z4�|�N����sy�	]�3����w~�������.�o���_ܙ�~8�Hv/J/�+��o���2���^��
?�m�re��Y��U|�����j��]U>O���<�ň��{s�k�����/چ��[9&q�\�U�L�>�^��G+�cS���q��������#�����y���]���]�T��Ӧ�ߵ����k��[]GC�>�>"�sz�����;m�V�s:U;9�>���w��}߷��h��y�q8�|�E�g^�k\��}C�)=_��X�<����rB�ͷ6Eq��z�sH�K�Ŧ��[�	�'��9e������}��x�>�:�=��~����!�Ce�g[].�(>Q��g�ulj���3���'��5^Nۣ���wY}����x����$�S/��^�M2�����?�����>a��|/�/_G#7��D媞�T���>��_����3r�->��"G�����8�}_��{L�Gk�+��p��ڧI�־�]M7������Kq��1�C�~��!���%��jp���;5n��	�x�?��?A˔8������H#���1�1�z_�������|���U��;�[V�d�;\��Y}׳j�h}����g�;[W���~j��W������������m�YOm�O
���>4���g3�c0O�������
"��:e�x9�g@߽s��Z9�Ի���p}���a�^�?B�W~$�����9��c���"r���^��b��=ڿ��*����n^����7�bw��ۑ����_����e�ߩv�9|�y~����U�� brŰ�=՞�u��?/�����6^���~գٺu�s�:�t��1�W��	]~@���>.��>��g�MiMirc�<S�Ր��7�{2M/���7I�s�V��G���������E�,.������+��?����{S��_��U}���u�D�?�?�Y���?������ܤ���b���g�+�7m���~�-�~a��}&��||j���'�ҏ�J�a��c\�3������������*މp�s5��w�\zH��N�I/�A�/xh��d����������X�sD~~�Z_\��`��x��b�O���{��s\.�\�l|��u��W���#��%�G>O��Ÿ��,����aw^C��~�W���U{�}��p�!�c�q�z�y�	{Fl���(g+?���e��E�+v�_S�{��gGn��^�W�1��1̭�b����4��o��}x����������������u(
���|������1���F�Ӯs�:�aw�<ΪZϺ�f�jW?����>zD�Ě@�	�_?Ú�/�����ml��,[�U��N��w��v��W�Q<:u��k����G:����A��V��J�T�U�a?��uu�&鈼��I�y����1�Y̋����&��^U��:�n*9U���p+���PPI*� ���H��hdPhApB�ATQPPm'p�vB��֦�v�m���F���o���������������o�}��{��Z{���W�g���z=��{[���#1䀭���7����/�Rѭ��?���)T�i�^mp�=���߽����A�Ƕx�VL��?�O��@��!p����^u���������d�x��y��S����8�R��R?�������t#��5�l���*NZ�g���n'�^��j��蹤�n'�u8����d�\eq{��uj��Q�ּݤ?k�����z7�ݲRU����C>Ǘt�;���!�T���}SǾ�%������J�'��<+>��+<|��hl�������=ԝ!֔����R����y�4�wƖz�7����g>�<r=2u�(L�ݫ{����#���A3����{ ��q���Ų~b���+����)�ٝ�!�/����j}���������f���s:�à�ƻ�p�����!�6S�㰜ip���H9_򾿝�;|K��/4T���7�"�I�2�ro��$��a����^�7ój_i�y�}�o^�{�����6���>��C?�T{��?���g�z��?��غ�p�|N;��#ǳa���B/ ��w'����^�E1��9s9���1���ys�m�CF�9�����.�{�O�'b�w�q�$�<�c,����<>�{;��sN���O���tr���k��j���%{�`X�
�y��D|�ٽ��?�ʮ;Q?�����Cdy��.�n�)�_?��o�Zof�:"�G�{���x�_���c�e��'w:Pa��W�>�^��������#��>��W����h�ǯ��U󸿷�;��(�����)�j��k{���>m��d��[�O���2w���ts���s;�)����vCB��1�Ú���={/��u��E���}.|���W��6|v��߈�X���[��oJ�{><d�oƠ+�>xY�ͭ�>ϦCp����~�����C�g`q�g��F������6���i����8��y���='������w��ܧZ}���xte'p���]{��a]�{\q�l�f�R�$5�9b۷���+zg�ߵ�\��?���]�~N�En�i|_��C�Kmݭ}Yc9�����|�wt�x����	�rR�<�{o�n���|!���ܙ]ܐ5�%p�%���|h,�gg��н��y7Ř�<��W��G�`�]�{�*}�R������rr����g^w�3�����ڌὪ��)qU�;A����_��V�2�_��c�w������]nΖ��Q�*?��+�y�^0��b�i,=�}��7��N��We'�� ���B�9�7==�5�}��	o�rc��ɟ�X���QԮ[����ý�<.pĭ SpWŝ��r}q���"����U�Ȳ+�r	{^��I���(���,���;�N2:(n�����l�k^��������o��=�8ב�CG���{?�S��Uv�a_@9�y$]�ep��rxf�e�����w����7��y,����r[l�g�/غ����ʉP�ٽ�f��h�9���b������"���漸��~��%�tt��}�©/�2��q���G��ۋbێt~P�k|T�Pn��{%���λ�ryB�;�����{�]r_��	P ��	�o��x����8�*�>�N�=b���T'�x��~�y�?�8W�,�_��~�
������$���!�]�o�O/��G�E���S�d�
�~u��cI}��(�1l�8�s����)��7�{6��윩�ӿmS��:���?�?P�a�ڟ��~����j^�y��,S��F��U����+�u����E�������0�oL�_�S�x q؀�8���Ώ���w��?S��,U�������?��w�y���j��>ذj��T�}]?C����Z%�-| ��8��:iOޟrOq�����xA�Ñ�'���=N����y	�X��-��޷��D�������}��'���np-���>�C�������� �4~��V��"8�7�ǯj��������I}��
��§�D��?Z}�&*�Ox�t�W��k#���կ���k�N�߁��^��h�nf'����{����[���_�eYގ��Z��=�B4O鐝�u�Y�-��^�e��
��+y����j��c\�Ģc�׽:�v���Y���]_�[�k��#���������Tz�}1��њ�Y�_���},�'�>Z����~��"hg��/�;x��!V	��y���u�?��B<_�c�����
W�zIF7�OH}�W�����ǩ��_�} �2��r\���{go��'��֬�u��W=��Ɗ������߻VU�ӓ������{z�SNd�$˷�jg���cӎ��0��y�����R����'��1M��_�O؆_!p�E�K�<ĸ ��U����?1��O��g������j���X\�5Y4��޹�y��:���!��%x�s�S�A���s�o�]��t�����L����Z�������%xܯ��.j��Ꮘ�f> �E��-��x���R��{k��3�1���G��P�g�.���o����;��r~�D1_����znw#���C9s�ӓ����KK�?S�'�˷���?n_[�[���^F�*�F��-�ul�}��#�����8#K���u��Q��K;�y��#�P�o�:�/��m�"?x~��=h�B�I�o��a��f����V�C��=ؔ��?�(�U��
���xAO�'���m�N���G5��ƥE�V�9�^�mE��1?Wq����{�خc��F�j�o�g��q�����ު��Ńf�mU�[�_�+��fhs6��{����J����W��v �?��+�ϭ;���}���������<
�syj���?a�>��s'�x���:%j;�^I}�U|E9�v��ԟ�?R��~�b1�W�-|���������*��x����Y*�k%��a��^�A����?r*S�<:�)�����7����T�.���X�1.�%����VэqX�5�<���ǳ�{!@���x��J��w����xm���bft���]���v�F���2��������U2��?�pS����\��Z�r��h[z�9����x�X\N��3�]܅��K�}��y!�v������E1�%��k�S�ll�
������L�g|{�)mo��xg������~:�r>6+�U���v�?oF�'�վ���{��n�3��@�]�K:Vy,�ת��rxC~#�$���ŵ�����{"��>޶�fmo<k�<;C�U�R��1���/ƛ�����4��_��g^C&�����K�����LNN��R_�\���b� ��9S���>��Z}��Tz��V ��� �B��;y]�m��&�v������z7�P��K��G�<�?_�an'�z�>w�����;:�L�7��c����(coN�?�97��OX}-��=<���q���*���:��g��w<ٹE�:�Y�~5���C�녊�����t_�����Mơ������y��c���w�@k��u����7�8_������OV:k}�/�潞��븲�>�}��a�_]��^`�C��K����~��������KD������n'ج�y�$γm�!��e�_e㽮n
�����g�A�L�UqX�Gh&Z��G���������M�#��y߳���ôO*�g5.��c:�y��{�[�&f�ck�2S���Tq"����N��H�U���1��4^��}��=�z��5OI�?��[S���b��_������+b�������r���XQ��7�g���P��Q�_���E?�>��L��t��?d�D�{xN�:OI�==���8�$x"r{����{��,�V�6G�>_�e�ߛ�g�3����qi�C1�O�M���g�7�O��j�M��s����1��MՃ���a��g��h������ ?"p�w8Ѽ5��c�/gǺ،E>�ap�$XK��y��>�ЄC� �yQ�O�f~-��b��-	�ʟPɟ�1Z�kX獖�?����\K����F��%���]^a߁���w|qA���{]�t�����C6䙟m��6�!������^��۽��,>�|��A�3�P���׻��`��{53<�'Y|�=U�Bρ�XKS�f�9�y~~�1����ҎA��/}C��j���W�?5��K�qX�c�y�LOE��(��)��ݮz�v��Q�G��gz��w����k�j�k���y�8r+u�^,x�������Tqבn�A>_��bQ{��1��?P�?�O�~�����Q痆���>q����,�G����M��xF�r��w
���j�R�I�U�y�/�/��w�A�9h�?&��Z�oih��3�߆x/��\�?�����un��3�ϲ8���`����ǵ���Y��u����'w��7�εq�n�v�q�jrdG���O�9?�'^0%?���l������-��.̎~�id=ξ�������j�_����C��b\��;�_�ۤߔ�w��5j��2>���U�'�\�k�V_��1�Ю���})���5.�y8܏�z鸎�g�uU������Gϋ)��{�Z�Y���H�h�����}Ю�Ͽ��_��v����_�q�ԯ��݄3�W���؟����/n��_h'�9������[�����!���n�]Z�{f�R�D~yR����t>g����/S~V�$Ï��Uu�Je?W�_���ϼ���	�0<Z��Oԏe~�� `�_�^��!����Uy&��m�L��+X���(��O�T�E��.�3<�	�����N��J���v����1{�\�>g�-�W9���sţ����\�k��7|	~��ߧ���+���e~��1^ו�T�����*:�|��@'��Ѥ~�_���=U��㹰?�b�R���>~�Ÿ2��T;vս��~�g���!�c��lv8�N�?jOrM>:�V�@��z����︁�	��tx����p]w���{���u��<1��ʟ�����A�y�Q�C�G��������h���3ƺ;��~��n,��nW<��w��ހC�M|j�b�X����D���O��f�����3b�W��>w��G�?ݿ��[�W��!����~^`�*n�E�y5�jG�\���G{]�R��Ծ��Ug{*��睑�h�oI���#�?z.U�J�o��Z��؊+���֔�y�=�����c�G��b?���*��� �|U�S&W��u�;� g���8�s���p��3�a��!��M	~�_���z���O;ت�]�����x0�$����x�8�>�)q�ey�
_�g��0�?ʩ1��W���U��1����ψm���qa/zs2.�kբ�μ�{�"rN��Ё�g|0�_��ʿZ�G��m�L�(�e���]ٷ�.����y�>qZ�|���0���߾�
g�.2x�C[�1�/�=��cj�0.yc���-1�=�g�'L~������>^��_%�+�����A3�w�"��s=��.b�����q>��_�}�E����?�k��1���E�Z��5�>����[�~�:bY�~=����!.�oE}�C?o����U����;_�}&ԯ��w~&�u������@��A*߲8�����t�xo����8��rX�C���L��[�G_�$��جn��y��.p��FΟ�1r�����W�`�#O����}̸�3�C����3�wU���!��'�:���?��Z��/��>��0o�թJͽR8�Ź�vg�<�;{a�{c�O?��>��6"�X�Z��4�5:l�'����Mȓg'힟�Gq�̉�]O��[��������^���q+~�:��)q�����a����%x��9՞������k]jp�E�ذ��>����.��f2�,���;>�o��Aț�ǈ�[}�%�G����6�{�ض�/��l�����ّ���{�3���no�@� -�8����`ҟ��c�%��E����-����+;�t�o�Ui}>W��>^�c�����}��������y��?/����c��ݱ�� �RZ���5���~���1�q�?6��a�*.F\~�R��*;�v�%���%.���S�7���&�x><��3%����s-���1�qo�.�^�g�?|j��#���S�{�#�ua�]�O��m����O�Wq:�/������g�3���W~ݍ�Z���y>��W�QcL�_���U���S?�E�@5/:��=�_�ϐ��?��_�,�����������ԝ�|^���4�	ț�������%^ɷ)�q��*�鸔����X~߾�ɗ�/.��^Ӻ��mm�>����3cL��b��c}}e,��Շ�^��Uz�M�S�Q�w.o�x�۷,����K��aG�������y�����_k}ǽ̈;�p��Ib\��R�վ�+)���I�����������'}yoq�ﴟ����1���1Z�����R��tZd�E�T�&����U�j_G�?A�M*O�k^������p�3�]g�bO�����On���x�f���^�~b<8� �ytR����'=���y���t�;cq��Ŵ��*��˥��s��G���G�9Gc�_�!���ψA��}��\��N��1�7�Xǃ�M�w�����ɇ��z��(�;?��R������w�"FL�Sb�Y�7����g�����1��k\��B��B}������ƻ
��'�s9|������)p�����1���׸%��53��/���Y�l�(������uM:(�����*��ʃ��˫�:U�gr��_�S�җ��.�5������]Z�X�"�S�����g�'�����������;q��ѷc�w�1n7z?�8y k�:��=��Z���^9Ǻ����^�)���V��~����:��Vr���?<Ft��/��YC.��H?�+h���z�ׂ�7r+�< ��~n��Յ��L�����O[���:Ւ��6�>�˽U�VvWe�y��'ʷg���Ԯ~L�C��$���o�0�o��w�#�^F�H���Ze��@���a*�-���<W�>e�D��p���=9u��b�0k�eO����7&�^ _����x�*�Eq+��bX'�{OR��E�������tp��Nu{@�|��ܬ>yC�	9rU���db_+9�v5����3��?[���� i���jW(2��y5<'�9Q=��UUAG�d�.��S\�.�c��t��o�~i��|9}�-�3{2�>�����/6<��\k�y�>��=̱����hgC���8�:��ޯ���ԸIf�y?+{�q��#�PT/@�C��-�����U�����~`��{-��z�F�
�)���F,��������8���Z�.��{D�1��W�3�>ό�<�Y&��R?GC>���-	����U��gu</�iruޟ������W���+?|����-�����|<�|!�-f~'�O�&�ysR�cs�����I��m�����hv������Tz^:�~��H�*x�f���|����	�1�ȩ�b�U�g���~~�������]�k��J��˃;�H��� /��QY|���<��'���c���'�����Y��|]_GJ�)�^��r���f��p?��&�aY����Y���}.j_eyA��*�G^��������W�1����U~z�Ҫ��<�^wv~`����GA����y�7��ۭ��^���H��i7�1��g|bl�QC�Beoc�~{�P�K��En���R�B�A����J��������������~���Q��!�'r=���hDڝ���m�nU�P�S�+�+�����
���Y�����g��Ԏ��`��XR?b������Z��UN��
{#�1x�c	ܿ�mN��+8�$�e����Т|��C���#�JYǕ�+��ap���1��}A�O��C^��!��E��y��j^��{R8�o�s����k?����_I����?N����n��S<د�z>���� ���_��~�_��_�ӷᳶVv��>�^y�I��������[֖���ͣ�i�e�>�Ôκ���պ���X_oe�89~~�~�*��t�x͙���q�3�9��_P�̻��o��77��W�5��JW���g�޲������g���e�N署�V�+�v^���)xԟ�z��/�q�������&���c�WЍ�<)���g����\!p�O�"�M��':޽y�����a�71��υ�H�x?�gG�ֳ
g���tv{��qw��jOFRg��|�;��]W�B�� �Ao�G��cil$�+?�֮�鸞���	���Uz����p^w,��эwo����-�����E�Ì�+��2>$�\쌱���?*�����[�3xV�Gc8�
��⪟��Ǭ��>c����,·��T��W�_�Çl������T9��*��m�z.�����>�꿞��쁈�>��.��~��	�$n�u�6�Ò�N�y�l�s^W$�Sc�/�=��>8{�C�-9����� �<?�-}L��7\���z�n���=��굛����{����ۼ<����oʋ��|?~Z�����|wu���3������H��g~R�g�9��|������c�!���;��ϴ��˷S�����-3nI��L*|sx�}����5�~n,��R=U�#ָ��5�Wۭ�9�����I�ߞ�z�T�?>d��k�� m��ܘ�'��r�/T�5{e�=|�[�C����E�y?�ڟ1g��|d��_�=��+�O�s{��������қ�7;C��z�����E�*,���w/�詰�<��sݗ)�@��m�{m��M���;i��"��9	�J�T��S��Z2���l7����tc|�p연��><����V�Y��*���=y����Y�����+~X��K�ŶU.�^w���,������]���`:X��G���5�m��WM��%��28K�a�ڭ�'��٧c�S}o���?{�˥U|^���ܮ�6�+���y1ް������Di����o|��g�O/���l��h����Ǥ���p�}*��7F�C�7�g��W���"�?����<[�/>��8��0�j�G�pfD�ؘ���u���G�����X/S�x�:���e�N�_��l߷����908	]�~��������}�;؉��=g1�3���OO�]���8����W��:yM����;�:�����b��
�+�6���E�A.�F�����\UF�]1�C�7�u�󿘗�:�������OT�����xa��gM�ˉ�5��~�կ�'
��q6.��վfY?3x��X���I�9������ψ�_Z�W+����|�)�bX�������B���9��؈1?���ۙ�Nϓ��#&����q'�V,ޟ���t�����k]�T�˾��x���s��,�P�#����'�?5��v}�U�����y?$�d�p����֝��ԇ���O��_y��~`�� '�~���g�!��+�5�)S<\���x����nN��1��]��(��q��w?!/�E1�e���B8��6�?���ڸQ��Ё�[��*���et�ǐ+��m��Ϗk|��	��1�w�t���9I}כн����Z�'ƶ���<���n��!�������z?y<��O���_S����A˫�x}����,�o�o�ra�8�^bq�D�1�e�m�c����I�v�z���X�s�'g��̱��_��F�lu��v��/C��|�sH+�����?ު��Mߧ��z�Ͽ���M��;�F�O~��O��1�ך���r�&��\��E~�.�?�����鰇Dn�x]eG�����^���8Ȧ��t��?x��S�ua���'x?7�su/��Q�>��@�d9h�w��Qoo�K��j�*���#@���g�H�����&tX�����p�yEO�{M�õ]�+��k��*O��M����J|y�H���������S7�����3�o�}u������C��������[��тՎҢy��w�3�v���}B?_"p=�xX����ܜϗ��7�ñf�kϳ��7�s�X�ǯr`�ܲ������xӲsL��8^��u�	��_����}\{�,���WW�xU~������B��t�˚���sV�C�����������c�O�����_�}w�O{���	<z���E��y?dp�w���սv>�;�q+�+���z/��_����?�?�68�+�t��c<���Da��b��{%tL����jU��|<�)��n��1��^�������0W寫��M��=����5.�x�8����G_0�{��>�;���~N��v١	��s1*7X\�<�?�{dR�}��D�����'d���k���}~�������d�N��ҿ��g�
	�#��"���c���� �b���d�ռ8������	������~s����|f�<��������l���ޠN�v���D�MϮ}���g��}P�3b�k�� �@��%�:��P�}��e�y��{��G�C��m	�e�j�f��
��W�VY}_��g����_΃�`!7���E�r:�ܓ����_��@�3��3�2�����悔c�����T��c�O3��c?Ў�I��3c<_�mǟ��a!�c6}����w6�x��oE�C�'����)�WƢ���Q����.��w���`J�k��zπ���ZS�UU����[:�Kc�.�~���Ӂ����!].�v�ǈ��?�y2{o���������?��sU��&C�ۚ���I?]n|0�|���o9�9\�5����N�����;�����{�G�g������Y�w��1���?��ڌ�}א�w�~��t��/h��{���O��y�����:�����+
<~���zy��g�`�$t`��'�}yl�I�>@����N�i�$T�j�
�������)�ޭ1ޏ�no�\�,�Ý�Q���xr{B��/k7��&�����'��<��nϬ�s�G��_��S�H�M���񽸅,�C�~Ǹ+��<�͎�H,�/�.p�>�'�;��dvW6^}�Ŕ8d8�(�ԽU���������k=�/�x�����ӟ��G���p��ξ�	Ǿ������S>y}�J��;����������mZ�ھ���=�|��'Q �η������z����1���~s���q�8��~eW��/�-�s����3�C�yS���������J�+�G�q7c�o3��w��~_�/���+y�џMo� �:�l��	��܁�'�v��X價�e���w��;;���G�O��N�3�&Ã|*�������Z���?���	���|]����?h��#�nx^�������W�z�b8��j�V�����>���Lo��~I�51?7%��|��6V�t�u��v�7ټ��y�/8���K�p��FQ���������jY��˓�{������e�w����+�
�E��_W{c��U�zs��y���w�xo�o���}���$���{�)׀?{�����p�lo)��V~�K~P��y[�S��k��{=�A�G�s�7�x^�w�ipm78�t�������q
�9�.=����>L���ߋ�z�����v�7a\��<p��u~f�t�g��v�8�ѹ^���'���s:L���pN�.�<�Y����g�eپ5[G����[�nݹ���G<U��k���#�y�V��.�b\��|�`��M�z��q�k<N�7��!��I��1R�1���X���O�|?���7?G�����A��Y��x.YR?��3uzW�����?�}��d���p�E�2�r.f�|ΗM�Ce�c���$�1/�~T<�R�I�p~��L?����������<�
:��)_i�|��I}�63;J�Iz��,^|I��-�^����?��ב���1��(I��������G,�ש�+�%(��+����a�;p$��.�<��3U����n������B�����ly�?�_�szܐ�M�B8b
�ϊ�~c�#��8��S/�W�O������t�<�nXJ�{�sb<�սX<���_#��zm|��Q���7�?��B�J�E\�����[}�oh���+��{3�~q���D��#����=އ~bΠ��<p��r����G��W�/�@v���迧.t����y����D]w�?d������a�<����p��΋�=�·���:���[=��=b1�L�?����+:�p��8Ǐ����3��v��^2����x!����.U>�8��3����+�g�}���׵�OH�ӊ�.ǘ���+��g~��b�i5�=�.�S�޷g�b����?�|Y1^�ۉ�9��c�~�j�_ݧ�y_�&x��O��vO<.p�EߋA�/ˇ�v�c��C�?�����c1̻�����ߩ���'��J�M��E�)��>���x���+����
����h>��*�au��{� wC����o/4���(����_�w������X|��S�S���~W%oy�����\'��N�s�鿿!�|��q��:������V�X:�.��''���������YO�����}B��	�'��[�'��������#r����o��!�%x*�󉞃P������ʇ���/��q��E�`E��b�{𽂫�u�o�;�]�E��k�C��'���\�T�!��U�+9��Ǻ�s��?�|ocծ�Px�?�S�k�z>�"��?�~U��Ew�D<wX����U���=1��J����^��:^�g΋\n�OW�K��ן��Yev�ɑ��ݼ]����~v�#d�c��;��/��U�b�?O�G������|=w&�\�tl���S��v���e�b�C�#�>�w3��4���Ƙ(���bk������yϷ���J��ո8~�?*�T�T��58�ZA��w��q�����9#����ݣ7#Ϸ�X�a*7�����hw�ߒx0n��lT9�ؾ��⤟�^��1U�v�/XxϪv+�"��v�#z}�iU�e¾c��Iإ��{�W�s|_�j\ap-����r�z��a*�v�<�x���I�}�����y�*'#��|U��=i��G�j^��U�b<	�Sח��u�r����w}��ܗ8=����ax*��������a��c�N�w�6\��}TnO�Ӯ�0��po�W�:�U����{ I�y�����֠?�;Hg|��������~��E}��8�>wZ}��o�8?qb�>��Q�H����Sx�g����/`�}1�')7���vžX��<���^xo�1�'����X�ځ,��_:Ə�j�!v�������-��m�0�7$x����c�
\��q]��ݓN�����F�#���O�[�+���;З�k��f�H�/�����u{���(�7^�������������C��]��g�?��O�p�CN��<���F��{��&��~Tŏ�x��@mTݧ�|U���
����}���z_5���vHf���3;�{����WyK����R?�g~!�F���%��o�xt��З������eq;��}�؃f�X��~Zl��L��t��ض����l#���t���vך����U�����~<ֿ{���������Ę�z��������V�H�{<�zaw���t_��;��D~?a^׃W
����S�#��Y�<�Sn�<�35.F��� ��h����-{9��N�|��C������6��¡�4VϹh��{ظO�i���^�L���^�	1�U~�ڱ
�������V~{E��w���}�����fQ�������Xw�J��aq�����������'��]�c��O��ײj\�/���Y,�4Ou��O�i����<U?U.dx��C����ϴ����#�ϻ�||:;���}⍆�㿏�����Cż�*>5u�����+�����1�?�!��?uO�Ez����r+?��������'���=����7��Cȝ3c��z����|��͗���1�����g�������'bQ�U�[���������=�I��[��9��C��"�cPFd�U�'] �<�U�t�
��h|'����>>�����Q�G�gU_�qj_U�����O�$��GbЧ�/��6�ߌ���;t�>����S���Y��*���ײ<����m�oz�1�d�K���óڿ?Ù@׿���ϲ{<���z�cx����+{�h,�)����ɸ��_��.��c��{to��y�*����<���R���������̌{J�ϰT~l��������0��߀�>�l�!�68�
�e�
�_�Ë~�S�� N7�!�#N�S�#?oX��Jg�����?*7�}���&l��V�{��{^C|���o��}@L���Q�w���ÚǼe�P*���� ��������W�<�����7Ȅ?�!'���������g�C�?�0��I}��*���]���	��Q��c׿��N�m��+����25d���ϟ��Wĉ����?�q��G��n�:S��	¹o��?"?\�{���$��)��-��*<����c�}��ݔ��#��P������|Z��?�����J�I-{߁�����`�i����_���Z�����<����߯�����:&�����.���X�w�#�ݔ�I�?�o�X��_��|��W���M�	��oeG�Av�c�����o��+ڟ����A}\Nj�2��oȤ*O���ƗW�A�ݪ��?g��j���������Ύ�l�O	��Ӳ���c�[���~� ��y�����J7�is~�w�����U>�ޢ�ޢ��Әg����~���$˗�~-��Uq����*gZ����9�g$��߫�Z��y^�sj�W������3{��Z���S�_�ϋ���:~��u�����T�RT����}�<�c���.�'=��?����Aٰ�����p������=l���
'x^�-����[��wck�1���n�w|��w��zCC������,�o�{��68����r���	��0V�G�Z}����˥;b�%�&���i��P=u"��*O����O�?p��������*��x���S��łW���������T�6{w���I�����<��_����yaq�Vէ������Ϥ��_to���X��˫���ʿ��2^�)��Y�����ɔG�*�W�u��qX�~k�z+�>�cս.,�c}�U��j?+�Q��i�yN�?��}{,��i�߳����'o��l$��qA��̐�cI7]�*���*ǲ<1�'��}k�<�{�����c��[w(���]�f�U�2鿯#�E�[���s{�2�2{8��]�����E�s�����4�wJ�@�׾f�m�����Ƙ��w�O����K���5�����֓�$��2�7Uߟ��U�)|վ�}�
w��5�r��C�ڙzo��<���F��N�c�^ъO����a�j>���NOmC��A�=�=��j_�y�����:��~����λ���P�۽b����Ġ�4OO�_�T�x�??:����I9ԟ_e�a�oW�3�Y^�籿�}B_���Z�G;��#��WS=X��r�ڧ������>s��1�\ov��İ_��)�"�c��:4_]�������O�?��F�_C�������"���׭y>P�G���A�窝L��������7^�!/�����|?us�K�+�/З#�T���y*���	�_��O���^S���|���롢%���'����6�W��!�vo��l�U�û4!7�!pƩ�k���|�ö�>g��*i���j?Hy[݇��o��\�����N�i�V�Hؙ����Z}��F-?�>钽gu��������X������ߧW݋�tS8�'��U�O���ގ�I�}S<��>�B�ϸԱ�]��f��)1��U��w�1�/������w~^����tf�ܾ�=s��K>z�qi���'���;���g�X}����l�#1ޏk�֝�/�o|}��3��[�gov?��9w���d�7�]:U^��H;�Q1-��S��[��ݩ�u���7ګ<��7�5�^i{��I}�7�3g\����^姊X�K�c'�9�_�g,���W���_]��|<�5����噽����������=r~�~2����~�LnO�C�_�=D����Q�*=���G��a����U�e�<Q��|6|���(�+��@�^�W���[�g�1�Q7�� |#�8��w�cn�q>���W�E��F�s�j�E,���d�3ܺW������lu���X;��㤋�W��b��E��~:;rykv���z���y�?+�xx�1x��c{9JS�3;;�]1�� O��a������ݏT~�(��~$�c+}3<N�#r�Q�+���+�C���{�^�w��:/m�1g���ǘ��S�z�0��\�0?��X�ψ���Z��H����w��r���H网��ev�}:���?A�=G���1<�y��?�������[As�J@���"?��T�^��<��V}����a�����vݾB�~���vV�Y�T
/�����9�?�>�"���v�������B����?Y�+���'���7��Z��Q���+<W��E������0szL������;~Q��3<��~�Kb�����خ��S��>+��kV�e�2�6VƟJ���y\��M�����׶j8�����W����/���[�'?W~wo���G<���7������<ժ�ٱ�N!�s*����}	~��ʞ'�O�����a�e��׼�O��E�w�8n��aߧ���b�#�N��~���{a#�z�z��{��*��Y��u=2���W������K�Wq�=1m�+\�e_=�\���A�}Q�*��_�1�O�{����
8�����b[�\%p����N��xo�Gc8��j���_c>?��|ߑ���������W}�{ԡ�d��蟙�q��-0�ϷŐ��3"�O�Em�GQ_�{\p�����ﷵ�?8�L��Gt�t�~���u��
����n��{+�x��E���0���u����������~�Ol�f����z*���d���2���<{B�W��G�؎"ݜ����~x���������-���1������M�5���<����9E��O�Ϸ���{]�Fݾ����2կ�}��ʷ����,����
O��x�>F���W�V���=?c~�+��卸���7���S?� ӟ��N��U�ϗ�m0O���C�k�3>��c5/�o�g]������V����J_W�Z"gR��B97j;!�sR��'�c|꯻WF]�z�E�	ם�Ig߯�Ը�*����\�G�{r��H�~��х��O�c��q�9�	��N�G�zp�>����=rn'T�SƓ���x=�p}�������&��Q��q�[c�۹,������{�nL���A��Z���������_��������6U�\���X��:��߻^�T�w��V���ݖ��h�ojM�*r~�v�߈�a���5U�M�P��9��qep�g�?��`p�C���v��?���}on�����u���8W۷��ƿ���}Z��1�6ծp��=3*7�Z؊�CN�]G��qU-������F��_8����з��~n�����X����ut�ԝ�G=�[��o�}tkm�k��>�P�`B;?{alݹ���W!�Z����?٦b#i��y�����<�����([�Og��^�w������q0��g}�[��}l�J̴?� ��]�]�>;�? r����l����R���]5;����P��?����O�g�F��e�~l���_����c|/1�
���7�?\'_;����<���go��=0���S�^���E�WRS��_�O��h�"~���g_�~��M�}2��3�|�yw�C?��{��zS��Y^(��u�qy�"��?b9)�~K�W'����s��>�����Ĺk��3���m������Was"�	]q�������.���Լ���N��|9����Ū�׳��>�k������#�S�n��,��񃞟����Iv�x��������g�����+?p���yҮ��}=e��_��:O=5��Lof��ߵ���V��'p�3�3�qO58�8X�����q&D�e���Y<��e�3{��C|�'[ �ׇ
����=���rI�� 1'����}f�OQ7{����_}���sʕ���\��K�nw�v��g���Vo�8�����7�%xP�����j=Rz��mlFnϻ~��G,�H��3橾������d��˥�1�CV�T�S�xY*�����8KO�ܮ�W,��;{��q]���Y<�����}$��W�D�W�9��԰A��s�M���t��|iB��~>���}�����i�ԣ�����}^����}�gG�zp��۟Z��;�Ku��������N���]?��U�5�Dx����</�W���E����}H�����GN����p�uU�Y�NP�<�N�_�mkk�/	~��]=�����oC~z@�������_�B�:鶤�,jgF,�-�kntxx�_�}��>��y),�{����oK�W|N��������o�~6�~?��o���1����>ώ?�g�ڥ���| �;��yX_����ʟ�������A��N�O��w�h^��n o�E��3�k?�/��=*p��f����:�]F7��~���ɸ*9���KE}�o a���gȱF�����7�cv?��A����]������݈����h��0�=2�5���\��rn��U�c�';�>�ZwN��w�?a���'��E���?m�?/�o�j⭭��M�?�iG8�(���^5�A_Ň�K>-��k��N����T�[oW�{���.g8.��hQz���h�Q8��X���z~Z�����Vr��>�y��An�
�C/Lڭ�pe7z��p��_�ȟ5�a�&���٩���i���3l���~�@·���?�E�gt]O/�x���l^�Q��}gٸ�?��p鸠W�szQ��Uy,^��::F��o���3b��'�S�R�zQ���)~��]�Yb��4����kԅ���q�z}�;�g�ɲ{��~��5UW�%��ף�{El��]�����=��<"�䦁����|~l�#f�U༗|��q���~�A�ԻXGj'+�T��L����:�>N�����_r�~ΒvC�/�}|���s��-}~U�z��&W�]Xw�a��xu�����Wk���G�q�ן�U~x����C_�{�m��er����1��G�7<�[��x��/8�1�>I�����>��Q<�ci���^̣�?�p���1��)��B��]��?x%��y�Z`.�fҮ���_��k�+�'��.��p9_�Y�g�{��7�3���lt��������r^�?r�P����a�������ߓg+	g�奆��ZUގ�kڽ�D��U������_~�〽�q΋�I8.�Kd9��Y�3�>/�����g?7��|��c��^#͗��`u�z}\ϑ֥&�v���Y����o�~����qP�y>!��!ȹ�M�����Ǣ?�O��`�G������g[��M���TN�^���=9�A�?l��G����f�=�ֻh~�5s[�O�۳T�_�'��h�(�+~�/�����{+������:½����o)�������>���oM6�	w���{B?�ҟ�O�>�����_���W�#汹ܫ��ٰ~�J����K�������ib��B�����!gDί5>��lrhM�l{
<���F�������Y\�S�����9��?q�Zm.f��{��W�~?����U�Vz�H�������ӪvY��	>u����9}�F�y�U����y�����w=��wM[�m���i)'��8�������T�����昶?�ƫ��
_�O3<�3<,�c�~$���eq|o�@v}���b����,��l~�������L,�ߓ�s�gĘ�Ys��*��b+�u�q�J��߈�]���}����.j�����l������bq�wD�W���1/��y�~zN��_e�y��W��>���>���B��;�?��������\�����W���=�<��~�}�}�����O��P����/O���<"W~v<V�K%}\���� �=�,�?Wy�xn���{��oA�+{�$p�ng>8���ċ(s���p�ڿ�/k����yAU^}���2���c��^���ِ�I�+�+�iG�q\��IطS��˒�}� ���+?��,�������;��9�¿��,��Ȫ}M���.h_�g�u]g��Y����/'�x��f�-;�(��K����}�yw�zD�4֤���W���Uz��i]�����K�_���	x��~��f�8�ڕ��/���l\/��w����^��ә�F?Ͼ��}����J�g��v �{����w3�ơ��Ϫ�'��,��cx���k^������4��[��S��:�*V�i����鲼�×u<չHţz��E���+�<��O�U����t��=����,;cl?Pnl�x^��{���Q�#O�A���Dye�Ϫ�Q��}��<�i6��{�P{2ލ�j�a/�x�E�ͯ�d��F�������о���a�=W��7!����?����<��J������U��S��W����7�!������|NӏkOk��꾻M��c�?+��,o��_�m��r����������0�չ�J?�K#ſ���>
�Oc+w��oJ�����ݟP�i�������,����T���ϭw.a\?���}D���'�Ufo8?����u�;|�~�r�?}wq�W��U�?89����f���Y����g�y�ᇏq��r}��,��4�݉�;�o6��an�#����j��?l�o��@�h}>W���4��̾�sp�_���ޛ=���,�hn�E~�u�uz<�z����)���}"���9|�w��3���=�����5�+�/����#��ҫs�S��a�M�[��M����<z}�o1�y,���}ߣ	��y��~���X�k���ʇ]����{�|�e~�*ޭ�:|n��z��n�����O�hGz=�$���n�1���]sA�乽c�C�V�ө��3W��*}�vi&=߃~�C1�'+��K�x7�v��?��;���� �q66��Ê?[�no��?�mt��uZu/(���ʮ��
݂|6�ϡ�_�Au~��}��5��<��E�wcǣ|N�~�UrR� J�L�'t^�*�}~����{EV�7�}4�Wu~�Z���3`N>_���h9�_Z�G�F���u=�{��?���>�L�z|�����o����~�}�r��>�3���q�tӹ[�� ���c9�25�@��?V�H=����`G�'�y��?���T�1�u��j�H\>.�_H�/��3����ݪ|��B\.ߚ�2�����n�,��Q\���\�oM����y'.���ָUu�z/LeG���c��1��?؀�8�qvL�#�_����.�ن�����Z���_H�T~��B����p���!�K�8������a���{4������qȷ�Z%��m\�������%Σ�1(���q�Gֻ2����k(>/ا��ֵ��<(��q��]݋�ZԞ���u�݅���u�O��!p�7?����ͦ�#>��~�ځ�Ƣ��؂�H_ߟ�П��!��>n�B>~e����/ p�-�O��V��l�p�1�p��@�	��_�9��_��oS��������/8�?_����P���z�����=0�EzN��f�0�����J���h�9��C��ړ�}�����|y��5�{ �񮂻���OX|\~�A��
9����>�ܴ�3Dn&�����}�~�_����j��U8>o�a-j\�꿮#�BF~w�k�x��	�^��|>'��ʶ}��O�����/�#����M�?�,�u��j���wk��J�U��j?�v2��A�C���b�[U�Z�Ϸ�O�A�"����?Y��Ͳ���R�/�ݓ�fI�˭���Uz���s���n�w����;��7�U�f��-�1�'�80v��K�����I�G�T��>&�?�|>���gx��z,�;��Ã���"ݼ�X��ɰ�9��Zwn'c��ucm}R�cV���a��΋1�����:(?T���v��Ý8���~��s~��I{����޽M�_�l�����~��EC��V��5ɸ��Q�u��oE�5�!|�*gX̏���R=2ċ�����w���O1�g�:�O�iyD���|dl�f�'p�W���}��OX�C�����6��2��:<������k��j��G��<�����8�{v�s��V����	�����?s��yq*7�8˖�����4��Z/�Ѽ�	qϭ|8����L�������cn5���Vt���|��W�p�perO�S���w�g�N�����b=���+�y����?��6����1ey&,����z�U�Kۭ���}5,���؍ʇ���*��	�)�l��u���|@���O�/��x�T}�^��}��������y�7���e��������p��o*�G��?�-�tf���H���"�w���E���^W�8ǋ5�|K>��I��V������]��o�<N��|�=��Ba�8���*<��}>�ÝoW�-]O�?Y���^���w1�qަ���1{�Ō��>�h��3��s������>*�f��n�a=~R�_��ixX\n��6�����"==��y���^kwJ��:'��{+zz�U����{���_�Kz�^���w��.��=֟���sj6���c���o���=�o�{�?��b�+�5���+c����yq?�IR_�����)�Y}�+��vE�Ǟ"�6���1>z�ß�=?���w�'k�ѺZ��$�O�^����g��*�"�s<��]p66��K@�w���Y��#>����Y�|�0������bZ%��֟����y�}���C�Cz�w��~�ʎ��^��y����'b�_�ч��c~b��\o>=���8�3ƻ!p� 6�%�})S�?5�$�#~>��~?O�'�n�\^��ӟ��|!��@�<��c>�~���?�龘ㅜP}A?6��G�J�ݎ�>��SΉP�,[�Z_��Z_aJ�6.�{~�٥���o�C�0~��_����H7緟ڝ!�^��ҾH��oj�o���֯ʯ��[�ޡѹ�*��3����~�(�+�߁~��To{;�Gn�4�z�v�ߗE��取�n�����c�)�\����i;��2{�ՏX�w���8l5�?l����)}jR���h��X뒇<�s�>��������7���ˎN��D�o�n�+�N����K,��ڭ�H3���y��,չo?��߻�����Oy�\/������;}�ӆޅ���Oh���O�S���f�G��T����S���Ý/_�>���V��et���nVW�����8�O\������b���G���1z�|��^;�s{9�kmo�������L���^7�e��j������ݪ��X+��������0u>�g���?��ZG����Fv_�����#��NU�M�W����o���N9����o���T���W������t]g�V��#&���'��?&�	��al�}�r�|����6�v����ex��q�=��!�
�#֊����Y�~�d��4�R����1�Wn�v�~0ƶ�Ӎ��>��<�z���Z���yV�k��a7���w׫Νi}��d��y�\�����6J=��*����L�W�+�t����E��a�x�E6�;cأ�*��8|f��վ&[G�����F���~	-Sڭ⿠�w��������������+�)~o��}���낿4.��dj��>���z�x+��Ǥ>�e�����c}I���0�w��)F|��Xѭ��CHg�:"p���o,���t&�^S�j�\������տ̫üM����O\�/�������;���)�Y���U<��vLC�G��������@�k~2�d��:�[���~S���:��G�7w8�+T��?��B^�/��j��J�!��d����Q������q�~�������ֻ�gώ�����~��m���_����B���np���_��>��U�}tu���Ǉc��*k���4^Ly���Kz�s���{h�w��������1��H�G���<��1ݴ��<��S������c��wU���g]�;����W���~ N���2{/��7η.��.���X��U����:ϫr[�_��WN׋;s�*��������o�F�zmn��m��1��Q���y��7�X������O�������C�ߠ:�^�/��ժ�2�u����(.�c�s��q��#(\�ou��q��W�{�%;������{��*�j]T~�ʏ�^�?�àW՞����x^�
�Cv���g����n�a�.�C����@���ٟ����xX���~�eپR��+aM�@�ߗ������Qy���y6�l���D�뼓..��˫e�����v:���kY��>H�w��d�a�a�Cv�=�3����m?�U�|!ʅ�*?��Ψ����)�0�[�x�5��O)��lq�{�{fo8~�Ni�K�gԃ����Q�<�JdrOi�pݣf���S���s��k��h��'�c���7��N����Y�iG�g&�]����~�=�*�y�������w�[C�+�W�#֘��dYvP���������:�׻˱Jh��>�B�{=��v `��7�3�����?�}J�="��X��py�������`��*����=��J?Vx"���|��U�5���� V�#?_��_6�]�9e��7���������}�+h��z��{��?��:��z]�~��|3���?��xA�[����:W��zϘ�]�>�O�F���W�L���(��o�~�N��4�}B}�=�k=��H��w���F#r}��e�����G���U�9���?�"��C{A倞Ϛ��Z��9�/�s�U�O�c�8�?��rq�Տ��QJ��?��v&��.�g� ��4�W��Ɲu݁�^֟5�t�ݲ,?���(�GGsy˼ӫm�7v8�����)�X��!�Á���Ǒ��ۃ=���o�}���;����Um��s�JOq���y�����Ln����*��*5~�rL���W�1�a����/��������*e|��I�0���:/�z
e97��I~Ѩh}�UA���we�Uyt�և����5�=5�y��/�C͓��B����� ��;�?�W{O�F���/���@;��/��Rωk\���=�v�w�δ]��bo����M�6��OX͗�W���:�1^ו]���kq�=K��7�7**�G��'�ؾ�:�^��x���~�cqW����\����
�����T�o�Og���N�m�W����{]�f�c۫��8�W=����Q�^�M�#VvnoS�T�.�`��e�W��H���I��9�����'~�(ذX���Φ~O���?穑ǩ�1�\�G	v��%���j��/�
עx _ `�=���g���X���W��uQ��*��*���K�:���O��q���w���+�j�u�~ ��ǵ;��WR_�-����78��5?S꫟꿴�@�������u��������,���)�>Ѣp���c|�"���?����c���zF��zߠ����e��=��3����J�L�<l�4���۫�r]�j=j�v�v������+��}� �� 0.M�e���� �\�a�ԿzBGa��H�������m�������w"_�,��*�1�6Ϗ�=B��P�{��������5�O���a�Af�h���99�k���8�W�a>���}���%p�#_����}�籰L��3����6��3���aO�lޙ懃Έ5�oo���\/�U�j���?�S��KG"��eq����G�_���c�|���2�w���W=��]ԟ!��K�]�������z������Q���v5)��Q�'�;e���k��@�����	�I�f8��5s4�~��ۅ������;���yW��B�;� �|β�;�c[����}�W%���������w�W���큦J�'�@G��+b���_ٟ��J���>��ڙ�?�c���C8'�v�]1��A��-��yg����u\���gz��_k1�˨�i��IP������U�B�^���O�V�����ϊ�<�n��,?��k8�J���g��_-�d�4μ(�t_�q�/�tF\��3Oz_%��<�O�����֍/o�ڞf��n�c�<�U���[5�J�g*���]/�����8���S����|8��Lǳ^��v�\�a�o~S,�-xA�0^A<P�S,n�T~T��������χ�T�D���1��s��W��S��O�Uv`�o�k��ǘ��_��>%�������6���X�o�h��|͗ ޯ�a�8�I�m����{�'��#�������:#5�r�����ߧ���ϴv��>�ϕ���}�<F���������O5�Ɵ3�4�m�s���[T�<��a��y"޹����{g�����p�k�1�?���Cg0�|D��\zz�=�V��mv�ؾ=��n���9�xw��=�Z2��p�O*���]�R_�T׽cQ�\ۼ��D?߸����d�Z[k�`��{$H������O�;�-���?_kv��?��-��^�}�+��mߤ�k���1�+����g�����yn�ks3S~cq����i.�u]�<D�y��3���C<��2����u���~o_䓋bLg���M��q�?��,^��V�+�6���w~��z�:���u~S������1���	��s��q;��o,{"?�?A?�οl����U�����sv����;�|�'A��#_�!��(�k��������#�_ڗ�}cq]�7���尷����_���cq��9S�}4ݽ�O�G���>N��g��e�yv������� x�\/�c<�\'��sO�yd�������<����ؗ�݅������1�W�v+��;�6c��iJ��ռ�����yA�a��7�@��W��Ӹϔ��Σβ̯����ذ4�����}�E�������:=例�h��Ӻ�����{s��q�|��'��L�3�A��>�}�����>�G08�̏����;�?��\Ϳ%ߢ�W�mT�ug�{uoS�S��� 7��q��9�l]���l��Җy�omC�-���5������J�%p�?G�V��i4N��wz�����2?�����qA>���տ�v��3�=6>�ȵۈa��[��<ٽ�}�������;�d������G�/:^�&ϭ�K�o���,>/���sc|?�������e��x)?=L�x0����o
����xُ�1�_S�U�T.������ݨ}��؂��	�0<�o�a�=jM�P?pE-:��c�q�qC�����*Ǹn�߃I�]_\���Ř��G�畞B����o��{���_�'�q�?E��~s��� ��88�>���R_�T��i������������7�� �/]'p�%�������}T8����ڠ�?��<i��V��~���NݺK"�_G��y�η�eqɈZ�����0,U�)�_fo8�W�(���K��f�|������ax>�?�6��C�3gqX���u��e�;������{A'�]7��׶��y:�#�z�f_�5�����y��f���*����諓q��/lPȒ�c���~Т��b��O����1~����~3�Qċ�(�����^��o���|���sF�z����U_�~��2�`�=�,��
 O��>n�/�����s��*�����u���^�;b|o!��o3��?�֙����r��=�K#��U�0�W�]U���_C�K]�/�x�<���Y��E�eq�ߝ��9߆Ͼ0�{$?�w<�Z�̣��[�_���0d�&����o��5�Q�qT�������r�a��R� �8[gJf����tS~V�\���tS�#:��_�����*?�����k�_Z|~_���~Vǁ����~(��<�U�0�]Q�W��(����龎�s"�����c��x�}2�7r�rR�y�߀|����p>{hkT�y����|c�/Ǟ�ϊG�~mo��g��Z2�29I�J.9��W��|m,�c��ș����=�ۣ;�g���[g���_v�����s���.�μ��������8�Ÿޕ�����5���7l\>�Y�,���3'��6ַ�W�u�d�"�߰�U�Î�=��GF�+}=����czn�b��o0ޫN=>=��h��6���G��l���^�ӽ��Y���˳�������a�>/��x^޺���Y�wζ�����/f�������S�e�:��߀t|d�-.�֬�|�,��N=�V�'��=Q�_/68׋�U/��czb����:��)�j���q������J��ݒ�q��E�������?V���?:���7�Ek��4N���z���s���u8�u���9���ҧ������:;��gc�?p����;;���ɸX���˛�����Un���-�	��cl��8�S���N��W\���	�����%����pE:��_�J�O͗��^�����yL�<���%x|\�/��E垮/�+�(���c9������/�E�=d�9��f�"���L>(\�n��u}
ޜ�����z��)�a�i^�'�������~y��G�,i���o������U>j��Ng�֣���Ɛ?����ٽ��ԸU$p�/�6�W�z�1�7�O��7� ����C��j��Z�CN��_-����l�n��h2^׃����Ͽ��V�陾��'���S"��[���`q~�<`�������S΅ql���k��>N��~?<��.����[�����N��V��l��'_�>�������5e���>��^�se��c�c��A���c|Ԏ�>[������>�)��L|�C^@�_��sVR��?�;b�B�!a�skW��j�i_2=�|�G��1�/����k�m+�����?������K�����ٝ�;�>jf�|��ӥn�Sy[�GV�����?q<�A�Ϡ��c�Ou�r_����ֿ�8����`g}c��e�y�ƛ�J��x)��V�[�;������ߊ�ʓl��������*���c���(�_�?�tq�]��t?'��������[�I�3����}B�¶��oX���ށ?�F��w:��������������[�ԝ=I��c�!�O�1(�������yzj�e�r>�0.~i�����-!�5�R���*^�d������Z�s>�v��O��A^#���J�����D.*yR�G�����\�3{o������g~ƴ��q�Mu^���Came~�#1��<d{U�C8|�л|�z������p�7����>1�A߀�X�O���?S�K{Z��}~m�>�qs�⼞o�V�A��f��i~�Cz}��գ�X2�r9P��,� �08��=��7�@��o�����1e��uW��
S�q�:��p��`�k��3[5�����	�R=��6r�ǭ1�w�8��>�Ur{-�u�*Ε�K���j�Ǹh}�;��k���G����oN����rA��O��������`?����k@�L��o�Anh� �˟��!��ߝԯ���{5+��؎��;������"pՃ�'�Ƶ*���/�C���u:T� �'d��{�+{[�3�>���of�������W�J�U�J�S�;�����~3�=��!�S�:������w	\�����ƫ��~^�W�qh>��)�3����;�����ZR��ey��*;����0��{yT�M��B��
���N��cl��_{����Gc|߬�)��J�����o~e!���m��6=����F6����}�Jθ�\�qڟ���a������X�G|n�Hs�=�K��t]Tr#bl���?�[�k�����1�S�� ��܆o�]Fύ-_�=��ǅ{�8�����?���m�A\��?ͣ���9�O�sTW��Ά����UE�H��.�C;-2;���&�̚�tr����Nm��^o3j��X�w�=o���K<��*g �q_��7U��m?2����w�f��A�W96E.ń���ɽb{���e��p�����dyP.�6����Sw�ה�_v/��~7�wb�_�߉X�c[��c�ߤ>�C�Tv�	��?���X����_�k��[�w�+_!p�)�+΢������������s��i|�g��n��h[�{����=�L����j��+�U����/+�O�W�%�۫b��g!���Ѻ����E_l����t��b�����c��y�H��ϋ}���s�����o�qq�]ŝ����;�맾����}B��������c�1�9��B��6��������/Řρz^��}(����ic��|-����W߯���)�X����vV����2��� F�rL�@��_38�0��>���8���gN�S�g�|H}������p��[��ٔ���;�@�剽o.��󅾽��W��U?�����&�|�	�	���wf9���K;�`�j|�%��1��δ��{�О����Oȳ�a�3}��Q�J����ɱ���͖�3�}����:�W�����a_u���<�?U?V���>��;�#:�|/��>1�̭s4z>���o��L�1�˶Ζ�>�~a_���t�����q�����Y���L]6e^ s�����O�75��� ����ϯ�E��]�~�C���S���*��s�g���ӆs�6�w�|2�*.F�Q�7���+�,��a����T�4?����f��D�@��d߭�?{i�2�t��q��z��I���`���l�g=�}$�\m���_ӏĜb�R����
�G��S�K�ݪ����m
>�� ��\��M��R�*��W��:o[�_���E?��G�i�n�����V �տ�8���4`��6�W	���;�tּϗF9/r��g��@���/��[�Ɨ	���S�*:`���5���},S����j��©Ή��=��ս����9����X��'S�Ο�����Q>���oe���^���+����&��T�)/tБX��~f��䀟�R<��>�|���G�wU>�<:]w���ן=�\�򿍭\���KclWlJ?%�u��X�ɾ��IZf�,�Y��䤾�[� �_���@�l���.Oher�m�<-�/W�AǛ�ϜX_�b
W�=ӳ��p�;��+y�Vu�z��w����lz�\�K7�wU���OE�l~+���K��I�^���P�u�5>���lxh_��z_���u�O��\s���?��_�Ё���u��?_c��>/���U�i�ͣ��5�����
t��wj7f����%i�D�o����jgN�װ8��������/�'�����6�����7Đ�sտ/p��.��uzBN��0�7�����1�����UY|]3�u$F����"���ץ]�>8��~��|O�M���w���\���h�k�'���5�V������2��&q^/��,�>��������,�����Y����շO��.�����O�������#�9z�?c~��5�~��W�D�Sǁ��Ƅ���D���4ԛ��|���7c���;:�~�뢺'����������EE*<,b|� ���r�f~����[�XR�����)��%�����J_8~�#�wO��+ݵ>�0z�5�h1��5�?\�Xt~������}�z��l28tb}�_��Z*�+�?'G��X�G�G�?��;��_lh�/p=W8�]~7�\���v�+�<�7]6{ol��g���;:L���pg>'pʁ��دE���W\�|�/p�wh�&[��0��Ox[�3|B���x�K�8����`�օ�#���"����ȷ�O�9[%7*8�<�E���|9\����_����t����[�zR?��.��ˈ;eyq�E,�to��������_lp<C�N����v���3�����3b8Gv���/�xh�N�v�8h��l|o��F�t:|E�|M�����1�?��>a��מ"p�[S�}k��9��V��R�yW�7���H�v:�?$��y���������^4�}�"���h�C�j�+��{����x�>��A>������#�pN|����}D���Mу(w&�ByC��b(^�c=#����x�E��~+�[f����͝7�������b��?��{��^W�״�N�~�������^���]���n�������7��k���%��n��>[�·�^2���zO4Kew�&�~Q�<q��g%7������or���H~.o-i7��:��^��?�H�;���g|�|V��m1�4=<ʣ��^�H���f1���O�����ZϾ��R�\vQ6��WgŸ����@����̬�'b���ي�g��\Rԯ��3�??|7���+H��F��8u�������fq=����X�p��)��]��*�~������v5�P�?�볶��?��riU\u�����j7���b_�����G����輜�,�U?��MۿWμ�?C?��t���;��y>�6�ʮF^�yJ�O�����F��G�x}�r�9���{qY��T?j���tS���1���4�;)��ޯ�^L�6��=�<�}�ޓ��ӂ�U�{��O�<%�?��}�O���mF�G�O�пC����2.�#�Ob,���Vه,n���X�w� �*^��Qd��gy��X���nǧ��ޘ)v>˲s|2�3�Ǜc��"�c�q}���*�5������7V������gY��K���1��,~���:.�n8�;xG�0+�Ga}΍1�9�2���3��k�,���e�ք�?k���W�~���	>!S\�7���ԧbx�d���^{N?��Y~�~O�x�3��<(���_|�o�v��7|o�櫿�a�#��g	��1�wWqX��'t�����"�_7ϧ:�>��k�v��DQ���<��i�|������3�r��H+�b��W����y�<�k��z��՟�������x�ꫯZ���]ol�g�g�#Y�����h�1��c�7�����A��������}٪���X���"|����x2^�y����r�L���t�-���MM�w�fǮ��Z�����P�Kz�2���}���'x�8x�w���z>��/�W�J��Y|$�gu���|��������=�|������ɳ��ܙ�k����<������^��cO��B_��K���sɇ�/��ï�E~��F;��V� پ�߭����q�?8�~E�Ӻ?ޟ/��T�M�_�>W�X��b�-��������?|�n@;ٽ�l��k$@�䏆���vWes!��<T1�{p0<_ܟ/����������L���(�{�u���cq~�/Z�AQ>C'�ߕ��u�vi�O���X%�??�˙������?؆Ͼf���#�����Ί�\b�ϰ��x9N��<|f~Eҟ���za�nFO�IU9��~(�qR�����y�r����G�Ϝ��=�����xo3���t�ʷ���!:����Z���#[�M������I}��6>Ú{U,λ���?8ߍ9���sXo��c�A~�z&�y����[�O�S�վ�~�=1>�C���sz�1����g����D�~9f՛�;Gb�Ժ������ض�����U�69�#��{UR��suY��#t ��ER����?�tf{.�J2{u������<>��g�6'Ё�ף�z��A���~�C������P�[c��V��N;��1�O���W�x���rO$.���Wѹ�߸�G�C�����?��pg�=��/�<�F�����j���!�d���؛I����'�~�]�~��c�x=��~/4�/����)��{K�]>{��H��H?��}���ӽ_*���+����i��T}~rK�Qj'dr���u�[�_����k}�7
nŌP�/N����G��w��\�)籿�+�S�˲v�}:���f������?q_ד����޹��W��j��3+~�<r:��K�Z�휪?������^��l`�],���q����A?�����o=������׌z�jP�����^xD��7��E��	�2��2��!�#�ym�/U�<�C����4��cGc��i���~�+�~����tߪ��y���k��t��Wz*�h�v$����U�ק,�ɧ%�?���߫���=/]���U�.緽����z~g��"���罯(ꇍ�j�P�a��t�?Ѽ �_��~]���}��q��z���)���|�yhO���ڟC�/��i~�gu��ڸڟ+r���״�c�7�鹪�t<������Wş,U~�S���������L�sU�"r�������G�\ �_����:p������C_�����K6^�+�k�=P��E�wt�����s�>�߿E}�u�|c���'�_�1"�8������MTv�<ո*~"��O�����?\U�+��^�՞��*پX�&�y>��N�p���/�o}h,�[W�1��X|�<3�A�<�-±gA��>zN��/W�����~a�^��cc;>���.��P;S��k�`ԏ��Ȳ������~P���t��㡼���{����ˑ?u~`֮�YЧ_���-���k����rf���/��z�c��k��\��x��m�m�����=�:�̟�����m��?���<u�U������h���������C1�KUk�����Tn@GC6a�5ފ~|��{$�C���k�d���d��2'������7�c;}x�x������g����)����N^&W#�;��*�G�퓬>����z_@ϧ	�vs��r=������tc=H��/�}��O>�~�}���v_}e?#_� �t4r~��?(����_N|W���E�F��1Q�{K?�7[7^:���|N,���՞���;k���^�uM~���U_WrR�m�>k�]�1��|����W��͛c�{�p�c �cx�g��m�b��챞�s1/�b�f�v�����lU��L�{�Ju���Wz�afo;~>gq.�y3���䳻�]䫵u8�} "��?�̿��2���s�;?�����>�~$��,�C�o�����y�\��V���U�X�K��+�\�s�n_F��wu<U�Zt�Ի��H�A�#������U�rLӏ�Y�C�����t������<Ṍ��@���M�~eN�ϋϣ�?�[�������+Y�]ϣ���apmS�P_{�����U8�s�M"GR��k���%�V|�v��[w~>֟?3�v��y��?_ո*i9u_O;u5?�����Y�[b��]r��^�UωE>yS��I?�nQ��,w	��א����~�;�窨��k^%g4�����gD������~i�+�:f�����+�Gn����cY�2G�K_��-z}̣�w��}}n,�E�:=���sO����cxo�[��#p�����~�)y�,n���z�������ޙ�1��~���O��H}���L:��{$���g�U�G�_U��Y��s���"?\`x��+�<�׏����k��[�m\*������x���*:T~u��>���t}������vW���/��:������<�;c�I�7�0�����K�[{_Ϭ�%'�DCsG�_H}����<�EQ�+��-�9�{<��O���;�sb�>G�1pv�\�6���������bi��*}�yw���6|�'��s�5�S�I��|�(꓎��gv���s�������= jW�=��ûL�c�A�?p�`s�y�C�ޞ멹�A�0.yf�rc��Q���U|��Uzrݹ>��V���1�����=�G�{��(�����d�~�Sc�ߦ�U��m(M����?W�e�Sᴿ��;�|N�[%�����c��k��ژ*��1���T��ӎp��28�r
�W���eq�Lΰ�>�ĕ՟oR���}ƾw��|���|]���]�3�tQ�������7����hw{�������G��N�J�T�|� �'�T[c��MWt@o�x��=����n�����&��3��vϏq^��wU��)����W*��82�	rz9;o��w����E֟0����<�N�U���b�n�vLc��g���U�+��o���*��}{�?W~H�Ϻ��]ҥ���V����oZ���h���-��Z�m?2C�C�gپ���Z,�#�9�X�t�T�J���%�g�1^�-�}��{��ϰ=��z���gq;M�a���G��Wz2�rXϻ!�����8샃}���x��E�z�F�q�������~n�&���J��\�M���k�����*<��Ǻ�-���"_b��C�"F��{���;��#���ot{��}�M���+R8���=V����u�*y�uU��)b<���0����=����.\+��:�?�P�k�J�i�/��b1o䒎G��l�ߒ���I%'+��{���\�O��ت�'p�ID�,b__����gޟ)s�59㸳އ���w������Y܇c|q���[���W ������f�\�Ϲ�s�nl�)�iOr~Y��.�<���k�[�ᵟ�E~�X�[n�_��޻��x��}����C���W�w�C��G��`�?F�������q����G�OU��H�U��^�?%���(y^��W��Ӽ��ӳ���gİN�����yL]/���.5[�	��q�u�#Zc�<e��2�_�x���>S�Yǥ~v��ҳ�?���@F���O���y)����ӑ����b,4��vlQ�,`?꽣�7�7�p����q�ޤ߳z��qb~�j_�����O���d�ֻ��/��*�}g������~_�{;*�za�:^ǣ��z����~g�.� �3^��r�WjvǬ�R�e����Ft~�t��藒�.�+���������&x����q��]��D�Xw��C1��>t�c����G��~f���N<~ޙ�ap�d�:�S�<��H�xͽ"��V~fo������o(�l6�l�������� ⢯��Y\�<ur,��������������U������I���U�V�&�3�ɻc���O�@K�������uծ���=����wv���������Z��*���]������>���x��g?]�T|����ˎ�������=:_X#��M�w(u]�;�z/��\ͻ����5U���$��߈q~��o�8��}��n�>�|E��v����9۸N�;��z���rf�=�81��S'�g���}7i����X�O���+_�ᰙT_7ݾ�����O�ߒ�e>>���3��(Ƶ��+������ܟ��<���s��c�[����j)�5��<��浝&������o��/��?���*�)��Ѧ�)��G�~"������3r�T>�c�v��S倖)~��>h����Au�/�Gб�w�M��@��������r�z\)�����?��GN�J���=V�{��3d��WvQ��@�Ӣ�KNg��������g�=��-��&��[צ����������m�&p�5t¡��7�rxU��C����N7�	��n÷|���H�_������c<kw5�l�k�{�ڙ*#t~iy>��ݩ�G��O^�y������uQ��~G�=ţ�W����p#U�9���c����S~s�K��J�k_�>\oE.W]Ϟ۶Ս�����+:���@�˻�_9���?\�_�3�~�<�(���?���/���߬�K�F�5�oc��M��4_�����+��|?�ƙ}��sN��E�⃾?�{q���T|��?��H���~
����������X���
�2{s3���uw��ԧ�u?3���Y�(/�{P#��#)�қU���_�<�K໋������T��X������oΪ����s4Y��i�:�OT�BOc��o�qCĐ���l�.������v�{.|~�>t+��H�Sb���5t�]�aX�����s@�����.����/�:O<��W�`kk��׻����%Y��q��6w3�h��ٔ��:.��^���ʟY?��1��^zTҮ㹠���~�j_@z5�w�_5^�y|\S� ����?�XW�[���GC�'Q��E׻�תvȞ^�s�}���vk�����c�����]�v����h�^�?����������>�En�z?g��������] �uU�_�Z_,�_p�����'�x����Or"�Y��p���'��t�X� �it�p�����~b��g*~m�����Y�E3�_ ��:}�!��3�u�y��w���L�{�*:k?���z���*��������������Sl���)_����~�z�譭�o�"?`.u]�\ͷڅ����t,��=��-����Z_�Nu~��[�S�����*D���.�ӎ�>�m�߹�B=���1��X*�W�����^c:0����d�~Y����h��S?%��c��~�.TN���`����������Y��= �_��G�'�O�o��xӔ�<������X䟰��oڟywb��$�Tvof�8���Z������v�ϮX�ﴺP�����.�)~$�g��y�����@����������}�꿪�S�I�r�\۲D�1������ò�(�]�i�?�E���:�ƥ���'��=]����G74�u���8�R^�_�;����=�z����KQ�W�T��*�)�}������y����������j�?����I�uk���՟@��e�g�_��[55�� �r������E~��;����!�����u���ϟ��{��X,��	������z����P�ܘ���ߧ���9�G������:��������A��;S�y��5_Q��:�@��9�p��)-��p�"��}���.�k}��S�<T�i����ҡ��U�1��q��cqާ����.���������*��8'��}}�>k���¯r@�վ�|r�<�����8����L690���K�~N������{����kj����g:ݎ�z�k��D��jgr<gƘ����|�m�َX���>�W���^�7ڇ��u��nu^��V��0xeN��,���	�l#��B^~A�O�onv8xJ�z,�?����QQ*�Д{�hϻ�~H�C/�<��%�?,��^��c�����I�sm��]���g'�}�^�״(���q�g%�ok��.�I����j�ڦ�+�e��"���|{�����O�O��F����X|�&ǐ�����`�����/�9��:��s sv���[`������J7��1�WO�a�}A�G��W�ֆo�E����wŘ�S���b�G����^�>���9X*?��ռ����{?�VďfOn��6��6����|�ywy�}�1փ���N�CA_�njg�|U~K������	���c?�^���s}�W�s���~N�W:���CBv�����U�Ю�~�Z�g��V���d���%'z�0����*��l��÷X�	�z(>���o�\��#��pl���C���qN��;c��Z�����������ǐ[����_�I�Ut�)uU_p�n7z�;��%�u��~~$���'���h�����=[WY���v&x ;���0�ϋE�>��W��:��?�1��Z�zF�g�������#~��O�q�ʾb�E� ��Џ��xuM��EQ�1��K�Ty?R{�����0��O%�.�k+�P�w��V�;:��w����i�xY���2�������>���}��������[����X����~���㪾�S���3�?�����ZS�õ��A��!�/J껼����)ϥ�w���dz��(�cS�K;���J�)x��|_������ v��-�T��8_�?�;��-I}����~c��׈���t���"�w���3��S���ɯ��K^���F����}���~�(η��W�kd\��#�y*ۏ���>�����Z���Q'�x��ƹ1���di�y!�J�T�1�`��y����{~��qW����~���S�)_Qn��{�g��`CH�ߵ���?�kx2�ּ��[y����E*�T~V��S��������<{�8d\[~dĦ��/c�Y}�?�h�������q�*~}]�����J-ڟ?�ñ�O�z�l�����[��`��c�A�yyC�Ñ�����j�����~��=��=$���(�+;d�|��soJ�p+��_o𬟕}K���?9T�gj��*�u���e�/�L�)���M��%�SU����*gt�R�7|D��y\ b�o�c���N�[gľ��Ÿ2:�|���վO��y�o�{�U�=�m��gUف��ï�WU<,�7U�Ka߭�����!_��=���������5ϙ��q�������3�:kx��r�����d��l?����|Ё�_����!^�-n����ﳸ�+���pa>���S��,n��>K�K}�����1����+;��N�u���*T~a�y<����G��<n��Fl����Y	�����/ǲL�(����ϗ�sT��p�L�VJ�)�����C�}�;���۝�C>"�����)��X���}m�b��"�Y�ߩ�o�n[a����u�s�>�U��o\��z?��K��?�y��rP��5�.���e�q8|�g��~f.�����q���᳟���o�.i�l�*?gǩ��{��C�/���?����c��4��q�8���ү����poW��Y~~e��b�|���o�C}_s��̯��"�"���-�0̙��k��H}^�:�q�T��S��Ce'��S�i��/�#�lp�?[�7������`���U��~��2��_�-����אO��|r�|F1^�+�vD�W����a~&>��U�m1�~�}��m8�b��cK���g�}
�1��ϔ/��V�̓���f2��p��1����꼳���N���a���{c�/~�W��T��e���� (J�Oc�}{�����:.�*��Z���dv��ᾴzo�!���4S9���Y������P�~"� 9��#~a,�>=~}�Y�Ϯ����"�su_�9V��$Ϋ����ئ��Ѣ����K�U����q�{�c��cؓ�I��9	�e������?z>]������uۮ��k֮��Y�ڟ��g���ŉ���t�Y���Zf� ���\�U��� ��_[��~\����>3����)L�s=�c��|�8�����t��]_G,��������̥���j�7��;�>�;�ѵ�۷��Zܯ�ѧ� �]���C`q<����Ջ}�֝��4�j���~�on��K��[�ҁ�c~�Q�V�����x�'�r����8��_c�j�U���v�>�'oĢ�!.���~���i�ov�y�o��h}���,������wR��Wlư����s���×�5������q��V�����xG���텭9�p����O�wꗦ�Q���_�c��~fWx<�um&o3y�����������5N�v ��������ѽޫ��l��O��cП����Qw�������-�v��ڜ�[,�i���k������)|�O��������Q�Z����<֟/�\��߀y�����6���9?T����g������ǰ޵��������	�dq�����N�����pQ���c���M���7��m5^��)��c����|�ʾe����O�C���7tܸ��X�����*>Kx�/�e��L���r.���:��O�\�M<���˔��	��F=��ɞooj��	~���dlˏ��D�gﻩ���;�V���S��{� 3Կ���1.�{o����Ͽ%p�1�˟��hkQ�W�����X+����N�ʎ��BV���2�y-{�N%�ݯ����^-���r��"��pRY��:T��`��6��14�a~=��߸<����c�ټg�J�N�?Q;L��ϲ��)r����_��K�=�~�F�#+}x?f��t`�c�3��9;���9ԟO������u�ߧ�<^�3�����֙��c��	��7�}�������\�{YvF�G�z�v<�e�_ݧL�q^�+����|���vo���~u����8�{fo�wbl��z\�-U������sbLO��Y1�ov����̣�aa?��I��G���/}[�l������*ϊ��.�����^���u��)�o�!���K�x�-w�am�?�P�i��e?���%\���0<�������~^�q�1�K���Eu�
�R�����|��w�!V���j�����:�X���ǚ����cq~!���4��a�������yQ���f~0֝j�y^�a~_�{Gb8�qy/�����7%��n�s�\�8�ϳ
^���c����ov��_��y�=�آ�ޮ��1I}��fw��w�4����ҿe�/A��#��3�����o����cL�Wϊ�o���/�F�����>�5�.��?��x~ig ��[衋b1?�@���@�wWl���n�u�x���~�S���cb|�9��&���ŉf�
kW�i�>�{��WĠomz��z�d�۩�#�O���f��ڲc!� g�U���]?j�s����8W>{k�����8���6�b����{�� ���z|��i�����7^��* �W���n��T����u3y��/K�U^Ӊ��]���{��-��!��:/��������^�t�h��`*�U���P<�V�X���@>@f�ǳ{��7���`g}V,��_�G�~~���6�<�?I�;=i�\�<s�[��3���o�֯����θ's�u$���xlcnp��w��F��ȷ��xx�_c{��a�^�~q�À�I�=~����h����Y|�Wy��Q8��߿��({O���g��Ԟ�z���
ݏ��o����R���H����E��C����7g�?���Vtc����b���{���4�{<*�U|����uwJ�֣�KW��m�}H����M6��z���	`��#�brO�V��|~=�����߇Ř߰��V�+p��ԸÔ|��OUy�S�!_��6��C��U�<>���ݳ��:�`2@�]���B�V~�,ϡ�{��aL�0:�������G��U��I��������}����(�	����L�S���w�ﾼ������;Dq��#��ou\�u��������~���7�0��<��y;�o�2U>����=��.���)y�#�T�aۄ��a�~1�A7�/�����u����Nڭ�;6��cݺ��3'����O��yǽ����x���3/��s����^P�U�6���w���z�).�9�^��/�ϐ�~?�o��~����->/چ��6���|��׏��~ T�n_GZ���1_�}��){t���¹.6�?�o�K߿��T<�~_A�j�N�׍?ְV�ǐ���J&g��������߷�"�]^U�V-����I����ݪ��}�q<�<�6�«�V�tޟ��ye������׫��I�����O��(��-;?������i*?��]�8��3���jok�T�T�n�_u;_�U��hL�g���}�cz��b�o����6oo�(�;{?^�| �A�B���6�kbx���s�=B,U��Ӎ����(ꯒ��h?ܓO{n�X~�����9��+���Ux��<��v$���2���Ҹ�;^腣I��7��:D�#�H}��j}��D���������7.�U/x����_����?=������ݙo��^�;t���T�nf?���%�#�}��,�^V_�W�����q�/;W��g����U�.ˇDٌ1�~T|���1��=�����l�=�W�쟏��������m ��o�m�CgQV����s|(�y_8���ӭ����r�G_��x���v|g�o�����g����{z���~�������g��}�h�?#�Cŷ(�����|d�t�����y�ũ?�sy��]}z{���c��4�~��~��W�6
8���6.�9��Tr���?���T�T����]_0���%x*�9���J~�?�f�|i�ҫ�~��;(��x�����3t?��8�i9�>վ��b`�'&�����r��x�����O���f�뺮�k��o�P�aj��%�-�y���6�_���~�}��b;Ww�=�v�gՃ�.[�BxnR���6.�g��>�Ӡf�\���y9�C6b��rYL8�r�4���Ԏcw��.���i�_��T��ޫ3�ΔcvOZIO�
���Gb���H�N&��1�'��>)�e��/O���2z3���xon��~���.p�]�����?O������>�y,΋�����gvN���rx�~硫��b(��`����/�==�v/d�u��?�i|��~��k��S:N�i����kx���Ku�</��O�;^[���T�`��U??۽1��u<����ǒ��bq~��h9?d�C��,·��҃{�s.�9I}����%*}W��&cfx�3�q�k�����C}�W	|w�aݨ�����Oi_	���Oİ����w�<�����\�������\�F�c�����ŐK���C�d��iQ�{K�Ikc�Ԏs��< 86b�Ͻ��g��r��7c,�('��ߥ���ử���>���?7��K�����k�}^b�)�u��0ȼ�
��1�b/�8�b�o���z3�㳾�W�9�n|E��<1-�>⌘g罾������	熲sd�=$ap�'�>��U?�~�r�K%ϗ�(\��U�E�T�]����c��޵d~�꼿��)�e
�y����=�����Vy�S�W�G��v��y������.���E�^9��vξ?����V���g�	J_��(L�E����z�.��xԯ�x>C�����S��*������%�+����0
�V�ʙ	�ߺ���M������5.�c�����{Th�;��O����w��ψ�K>9��s����#��a��"�Y�n���ηr�;5�T�K�~C8�ZB�n���f�y�@������O�w��I�3:j���d\a��9���'�!1�G��U1��[?�F�=߇�u��A�C�U��T=�z%�cz}�S�������G!xQ��C�+�'�g��!���P��bo�i1���Ƌ25�@��X5�Oj?Ü}��/���Y���������i����	h ���$<�_��7���v+8�Ƌy����Ӷ� ����U��zti^���T�S�ӧ�Me��2}��O��2<�߀�c�p���=zd�~K����7*{��gj>��_�/ĠW �4�\�_S�W���nz��墉���3��d����^����v����?%�9��X�+��=|~�vsܧ��|���|*�#ͧZ<�����?�m�j?�������sv���]1�=4����8Ϸ��nO����B�2X'���Q;���Ǜ���e�ep����W��u�|�~��E}λ��z��w�*곸_����h*7t}����}D�u���x\����A�gJ�o����\��8��b��x�K�������oW�빴����}�A�?��Q�/�~|�����E���r$�^�	��T��e��cQުL$g��=�J��r��3,'�/�����Sg~��+���~_f�(m"ށ�9���|	�Ụ�#*{{3�=7���X+�d|��2��}���dv�����;�?�˦����?�ƥtP<j]�����z�#������e/�F�S�|>��</sI,�_�g�e��>�ٽcL�U���v��(��"��+�� ���eW�%����~����=��#��B��K�l$�]nTvuqHyO�k�x�9��5��S��s}��Qg�x_��Qgtv<X�s���G9-����d�SN��y�,S�	,;cl�[��b˿=�|�����/��>�?x>�,�s���+�����9���Ye'�V����<K�[~=���/��R��}e,�ޗ�ɱ�>����9����K�_���)�P�#R~f?N7��s�>,\���k�j��X�|\R��U���~�ʏ}w� �7����?0�0/��}�a���?gq��R?��+���� �>d|e�y~�~���m�/��s��W�Y�.��X\N�f��͎���N7�?_�JS]�ψ��򔸶����x�g��'b�߰>���������e���8����EW�#��*nX�?xs��������p;��,.�;��~�؍���v�OX��Ý}�gL����{h�_�y��q1޿�}�Z����J=����w�?��2;��cV��ݾ�s�O��y��G�7�nW�	���1-^\�Ϻ��	�ɱ���j�2������ɬ�[��^��Igq~��~������׋���6\��~T=²�Ϝ����v��Ɋ�'�.��v�	������?���9bە�C�}��)��2���������G������r~����������{���=�G+	|g�r&�בE�F�@��P�<8��gN�kc�+�Ǖ��Q�e���I�=~���Ok�%7'���M�g~�;�r��ؾ������������5�o���z��}^��X�R�s:�������a�أ�1��r�}}U��_����>e��#���ۛ��������'�ȷ���K��3u�Z�e�}elݻ:;l�zҭ�G�}��W՟���r��3$�~I��}_����K0�
���A��!��vK�W�C�̏��/W��>Y|M��F��ծc�����g?��@�O�����*�����35O���v�~V�y,ίߧ��B�!����y(�N�Ι]�򰢃�������Ol�ف� �ݧ��}C��5nU���N�I�`_u\W&x`���^i�G���	�:��l�o�G�������V�v�ᭉ�H�L�����5����=�tf�=�����8i%���܁w)���{�����#�p[l�Jk����+��v~���\�W�ŧ�^���8�u]ѡ�/�c��k�����u��������e淡>�{B*;J�Wq"]_l����n2���˷#��yT�{�� �3o%?+=[����7�썖��l3�����5C8�8�=S�oQ8���x��@�c��V�k��wڀfO܆��5��e��q��o�?��T�N��#=���G;�~O��c�m����+�>��K��?�����rw�d�F<t����+���o�~'��j��ۼ|����������|�>����9	�D~^��{�������5��j�*����?��ý�H�8�y��z�@H=���>���3���ܮ��^�y��=���İw?Z��x
���g�'I���Ճ~(r�_�վ����0xE��]��.�k^�v�qO:�.��Ȭ��A����=O��O����˱�?��1�_��_=βW�k؟��W�������}��w߳����I�W� >O�����F���#�L��lp}�`f������X^Q]m�+:h��d�~!���A���Vt�o��V�B��m1�z�ϫ�{�S9�y=�������m�ʗ���x����+�+�x��1>w�y���:�o}�<�qg��3[�.�O�����́���`},�����S�������ƙ}���M	����؅�Ń�ȷ�/@�*|���i\~U���Y�7+<�7Z4���g���!��r��?��aOB_�"p��7Ű�_7��j���z��?�'{U����o�Xa��o�g@ϯ��>�b����2���'��_4��hr�5�H�e�
Ń����q����~�^ų�a��y�������3oZ������7ǰ�?���g\��w&�q>a�u������ʗZ��3��3s[	?g�k"�6��
�s*�b��l�����e����H�=	~�7�o���OTٝ�*O��~�+�b�(�4��{��^�5��p�{�X\������{�_��~6�u��G�:�R����
���_��߿�qn����q��C�>d���0ot����i��g<���df7R+�.�����|�?vxw�b?��xֱ��j}�7��w������Q賘���^F���~��}_���Uz�H~6�yv^��Q˔uT��(���d���������Z�3�[���ؿK���hp��a� O{���|R��U�S�O���Ǵ}��z=���ɸ�p_�����:z�:��/�B�_�HeVp_����^�>�����d��;�AW��L�P�������߯�O9�D�wTx*x��{'�w�o�ߌ{!�1��c�g�/T�T�k2}��U�|w�����W�}w�ӭ��q_9�V9��˵����/�+:���X�OU��������A��Ԏ�R����?�(?%p����_���p7�j�-��I?=N�|��j6�r
��8`�z�2��4�;�܌E:;_U�S-:.���"�+E�y��<����y�*l����B�gz��TyB<���{c���^�v��W���}D�O��N�c��U��������4���q?gW��z���3|�ͱ�3bGȇ|`��U��	�g�Ǳ�g]p?�g5�>���/�����|/*��z[ş�W��F�y��g��[�~�إ�_N��O��M���)����Sm�L�j��z����Ѓ�ך������t�A}�����w�p緞�}lǍu���w�!!ߥ�g��w�X2j=��\%ߪ����P��3=.�Oo����6�f�ܭ~�j�E����b����������P�Vף� �>��uYR?��ZG������/]/�z�g��u��c\'�X��|k|������T�!�{B���������Y,�7�NV<ڟ����x��/��s�����wS�E+�_��W=���g�8����>��K�;`����<�S������ԏ7��n&��D�?ap���C��|kW�eh}ŝ��q1��B�_��I.38�2=��{+~�q!�[���+�Y������
�_o�夦�v��S�J~�%�.r� ;��z��U��}}�6h�r�?!��{;m�ϰ���il����~���\��uu]�w�+Mѳ,G����^���O������B�a��*��ʓ��ҋ\3?_8��m�g�J�p��,��^����'���S휩�*�Pv?�^�'��\��A����uQ�ϔ�N�+;��'�T�98����C�Z��B��$�+�C�x+�\��y�Y�}�����S��g���8}�b[�L9/��{�~�!���8�M�X�;�[m�β��}?���|<�v��^��Q��?�o�j�`�7�*�}wN�_�c����N���*N��g�9�yL�sO9Iƹ�I1.^�sa�������������ݯ���������"h�O��#~Ϸa�u�����+���P��x���~C��O�ؽ?G"��{k��6���>�CR���{�2���M���ؾ�V�{m�N�`|���3bL�v셏'�}��c�1���u6.�b~�_1����S�H�3F.����~ׄ�?��M��=�Ѿ��>�F��K���7���0��}�(�o�0���^�aN�w�ǽH��z=/jE����/��.�,~�L?*���� ����K���x�y�WںC�/Sxe�T�W�`>ծ`>��u�<�y����^uKf�T�Y�o�g�;&����������)��1����6�y �c��������R/�9��ߣ��2ފ�,;"��G㧊�t��)�w���Ϡ�U�Wv��	���:��KB�[b���7���~��"�i�{|\��y"�<=�08�;���R�+9j�2~�y����0ȱʞ��B?a��Q��~l�'�N�O��N?��)Ur�����]1>G���r��T�Ou���e�JfO�:%߸�㼟c����`�y�E���5I?�<��E~&}�{�?�v<���c��������5_���B�����G��	t`������<�\�c"��|����G:��_�@����z!�+_������\��l����>_�����XN����W�w���!��]ʱ�c<�\׻�!��9�P��ȏ�I�C�CWa�j\i��v��3˯`�:|��ʻ[u�t~QR����1��޺^fQ�'��E��#���C��[g�_>�6��>�����tjL��X;8o���Gt]d�|�����h�_i�W�� ^�k�h�Ͼ�{_��w��ΝL~j}��U��,�����}��Lex��V�Q?s����Y� ��U��q]`�+z�.�������7�?y��!�i��+�9�[c�~d�CV龏���V�+� ���{b��h^���_k��H�������&�!������ֲT��U��*xe�S�|_�м�֯������D��a�U�d�,Nm��|V�3���7Dn'�^���PA��?��>�6�b�?��-~^F�x�U�+9o5��&��z��P��ߐ��W;��1�[���+�{ �8}\�߯�?3�|i�3���q��n������5;5�~N�CfO�^�q#��"���Բ}�T�K�ת�WqoW�A���{�~������x�H��|1`Y~�T��۩��Tp��x����.'������������t�-���!��I����>�u�{�.�S��|�[�Z���5�����W������굛c�?�6��"��U�]t?�3�m:�O}o�<��L}��UU�h?����>j�j]���Y?���T������F�8��^��bq�P�y�<��{:�O�ΐ��<�"+����x��u������T��:¾�a���O����a��s��������x?��#C������ͱȇz�ܚ�;b��ί�P�o�WƁ���a�up����.�'�.�\x��j�z�u쟇'���*�R�>X�J��*�?�p��=9*����S�C��v���2?LX�G��Z��X;o�!��~�~��?��t����#p���1������_��d^�z_�=���oe��4_��#��E8���}���=G��_�yX���}���/�)�}�<��8T��'p=������s�[A����@���'������~��ŭ���HA��ߦ�����Z�����z��|��z��ٴ��imϹ�^�k�V��l^K��@�T���E�
m�N��>Q�X+�W�s��������>��Z�z���8g�49��v>�n�X}�=���Kꦏv~q#��L�3�=��
8������U��_����;�[�o����?�G��:����F��j�_P>V~l��u�Gם�o��v �<?_�yU��]%�*�������?pJ�r�������z��~	�cv���=��Q�m������������7��A�r@�/�Ǳu~n��|E��"���;#緰~j���_Ģ��R_�3���M��c�?�W��,�G~�=~M?��]��CT9���w����6�_��_�?��	k?�~���+Ř���b}��W:���}�O�ts;����*i��z�l�s���
���V�k���W}�t���x^��십��l}e��;n�S����N�*�X�>{�q���&�[ǝs��ͽ�ő�_�H��3ȁ?j�mLk�?�������ύ�"ri�z��>��?�_���W��!i3�#L�/�T�g�<��1�+�4�1!u�^���l?�����{;g%�}�y0j�����ƚ�"?��xQ*y���D�)U\uj~E�՟�������3���O3�sJ?UoN����VE��_�}Y���Y�3��ϥ��m�}5��zn�Z׏�ϐ�cq�*�Z��dvc��L}M��Y�W��K���?����ύ�����<��^[��Ͳ����І��������������Q^˲<"է��V�%y>�!o����>|����_�ݿ�/O�%ў�w�>n��׮��w~!�?��=o����d�ψ1�p�����O���1�,ƥ��L�L����Ur���y�1w6�cվR�Wy,U>!�r�o��T��u^��1��P8���:������eٺP�̾[��+{�z�Fwp: o���b�g��5:��?�^�cG��k���7]�:����jOR.Ǯ>u_�Ў���)�b؏�C|l��Ѽ�̯R��#��m1�Gu?[�e�V���/�����\�}z}�!�7 ��!����b�nN�s�G�����q.��<�|��;e����7F}.�D��.��:c���ڊ���r�(�~���~k}����fO����������M��m��?m��{;q?��6��gT�~VqU�u*.�sV�A�Bv��zJ��=����S�nծ��+��t�ٿ���n��<�X��\��ߦ��Wx������z���P��pS&o��ކ��6CL��/n?�y�������W?g5^�+�F~/��y�ez0�cV_�g�����J^:�»K��J8_���}u96���c�:˯@��	|oǋ5�q��<��w���;҃*Ovm�e���=+��ҡʏ����Y����������"���J�������x_Vȱ�f+����ʍf�������{p����������g�u
���>���ԟj�C_c�B�>��ϒ���z<e��&��ǹ������,���Xa�e��:��{uZ����?���������/~@�y&Z_��Y�^ծ�+)��k1������o���ϣvr������������ڶ.g?"p��Q�S��3�?�����ۙO�����=ؕ���t����GݗN�_�8���,�s"���W8��d�?������.�^�/ݏ�ߕ��y��mL]G<�A��t��y5�j_�:^���"Y�}�ܣ;k{굶&gM^�<~���w��}(���'�g����ֻi������%�iO����p��c����Z��_f�h����_��k�c�<>�ׇ��	tC�p���&�q�Tx���r}��-��5�t��U~�2`V�}r:3��ɱj�����5	�|$���i��֝��(~/�&����矈�|��w���>���Ҏo�:�~~E����ʋ�����?�qi������Y�����>��ǫ�^��O�S{��k�E��0r���f�U?��1������ٟ�/�]��f�g���&�M��8?����x\k�u/h��ǝ��R<���o�G����ėW�IX}���;�{���E������9�����"��C_�-Y|a�կ�aP�
�􈶩�y�~�\�+�����X</Ӟ��לr��r�o�X��/x�[�������W�[���?0ծ�㵴j\:�!�.�F��RqW�����	*o��������T{/�o��T��qlj'��;���L���M��6�eOK��<;����O�AU�a�;��}J��،:|�[gt;��6���*����������>�q�#W�'{_Fg���r�����t8�d�e���;c,'�~���l�V���n4;p�1��~�<�����~�U;2�'�߫���~M�����]����Wu�Ƙ���An��CS��D���1b������<_�1�+n�8��j�B�v�����av�8�F�o[�O���J�_�q��_{]lŜ��;2����}�i����_u^��_�Yo�2�������#��\<�����U��rJ���~��p�0>�~�j�Y�U�[���v�wC��!����k`�C�`�sg,�?���[o{���ּ���u=ɷ�>��ynO�}�dﭮ�F���gp�'Q�C���=���:��o8߃�nx8��Ÿl��M���H�k�e퇥>�p�2�S���D��y|���m���S��y͛R����=`WƘoI���ٸ�J�Z�}
�|"������ۻ�|U�������ga���<U�W�ƶ�P>����y�� ��9�A���t`�%��]E����f�_/���M�?�'o�x��?6�?�Oݬ��h~��_~]�X���'��e��ӿ���C��wA�}�=�m����rR��+{W9Ԉ�}2i�D�$ap�[�e(�b;F��k�o�����E��)�z�?�>�}��y���J^�ꯢ��S#��"��=N�^�y�q��>�s�슱\zkl��Cg{U�����O�vu�dq�y�Z����X�[�[�q���G��ٺsgR���@�g!�4_�1�[����#Ur��[�e�����c���y�j�V���_���.cdȥ����JnT���W+L�t����~�����q>T��������ű8�į���}T�cv��q��1���Ц��#�j��}ON賌?�v������"��G-�_n���|X���q�×�3i���j�V��X*?g5.����X�G�}���x?i���9;|�����qW,��V�h>����!��>�������0
�[{_-��wE���W�~yΙu����>S���7��e�xdv���x�#��{�����q���k�>��6c|sf���mJ�9�1�ono�E�".�S�W|��{E>9�q�Ux*~[��1�2���w���ʃ����N�t���~��/W�O�c�W�F�_TЁ~\��z��?)���Ǹ�'�/�v����<���`�r,�~�fq=ru�޾#�V�;o�3�3����v]n�7Vٷ��Y�Ժ���tv�v)qN]_~�{e_��ߙ���,���yq��孺ҭ�+f�t�����:����Wtc����~��,�]Q����{�֯�g������������_���zO��Gf���]�M�Ϯ�E������.gV�	F����HǛ��_��;���5�s������}��gĠ���;�_�7����� l�`�k��b\rWχ*�j�
��#���X'���:2����G���_ޖ.�f���uļ�y�~B�7I�:9��>^ʁe�G���V��N����������J_`=�v����(�����݇��V�5��Ç�h����9�Q�Ε=������{y/�������������!��X���g&oq�qv�k�r�|���x=���+&��2��ϼ�����t>�Υj�Y���u�e�3����OL��lwY�I���W�ϑ�_��<F̣��ߙ=��ʳ"?���Ϫ���������;>�k�G񳸿��X`��]>7S���=#��c����ռ�7/`��߫�%*<j_M���:�#~�է~::����w�`�W,ί�I�7Ű�6�������P��<#r�̒��gI}ʵ��x?���q\#pʱe�d��n�<���u�����N�j�j}�Ü$n��~X����Cy��1μ5���1=��.����p*�����������s�~i����\N����������	���>����X�C�&�Q�d}O�X�g���]��<.pݿk}��W������:���vZ��#�O���~�L�*��~^f}�k����MeO旛�x^x��1^_ڮ��y��g�Ϝ o��攇�F��%E����k[�?�E���b?�/�����o|6����\mC�Y�w��*?
��o�_�}��uW��ir��؎�>_�������po��k���c�3W��`�W�_�P�!|@�7F���?jO>����]Gls|��oQ �*�|&/��L�7������yz��+~$�{��'�o�������U�%�[����;����v��޹߉:��P7y���Z�.�qq�6#�s�#��~��/�g�V>��B�w>��藮ӿm��?��֝W'��%;�����H껿zo���(���}�0�5�J6~ck~�#�_]����|���չ�����������)����fqy�{�f1��i?Uns�SG8�#?M���gE~�~6^��p��#:ȱ,h������c��2�W�ϋ�6!�����ɷ��q����������/�<�|x �\H�g�˺O����5&[���;��r8���_��<��E�{[��^�e0k��x��[���غ�q��+�7�d�<&��[���@�y�(�\u5۽4F��g��gfM�DM��@�_���?G���N���靖ܙ�?���.�K%��Y���� �}�������Q\����7i��/��_�����5������xD�߫��[%7��x,�!�O�vy.�����{"����|�J����c�.�[��?|���}�����?b|F����ЙX�H��v��y�-3u]�.օ�-��YV����U�}�x֝�X2=x$�}�N��W�J����}�N���C�䘞��_���,S�%��y����ǽ=��SG6^�#.��g1�����8^V���O?)t�k��ዂ�-��l���y���؎m���}J[���G���T���5l��!��AE�c͛b�l��/�������OR�+����yڏN�_�i+x�Gb<��~o_��<�����JuoF_&�3�������ڸE��SxEO��{z�C��:_:.� >�i��A����q��>��N�X?��^�ke*��_��O��y��٩[��5ǒ��?_�-�ߪ����v��_�f����y���؏�0�߳���]�����7�^*9�m�j�Ͼ_ca[����e�k�r�G��&�w����)����Y�����m�����)��=��}6[d�7&���x=>������~]��{1~������f��'�X�����U}�5�W����K�����:��GNٻc�A�M����'r���oS�;`o >y�՟%���kYO�O�<B�������G�ꩱ�KW��L��U������gG�}��:��	����}�v9Vɷ5�{�r ����<��V9���;�����]������q��%���g���;\���W�����I}�mS����i*�ٮ�w�h�S�"�'9�oV��gG�޵������`�B2��}CY��>�~��Յ	�3�>�����k���G�oU�V�o�pV���wq�׽����w~���8WE�����_�������8�.7���r#���7N�g?���}�~��D�`���y�W���P,λ�ũ��<ԹW�����>�t#�-�O-ۧg���er&�3h���A{s{u��7{]�מ"WON�Wr��W���y�,���z��,�︾�lp�j�$p��Wv��1�y���k1-�M�g��ǥu��x��W��v�:9�󻯏���q}y^���o�_����k�
�����x�¯E���yW���t�*�����1�̟�|K>���?��|�m�x��]5~��+�8����C�����?�5��ު/��$����;葝�͇%��������	��Q_c��*.�6V�a�=o�ء�ϫv���/iW�3%���7�S�c~���)[���C|C���CO�<�����]�o��Z�#m�����{���L�/��S���{3x����n��k��7���k��)��������=}���)�_�[����z]�{��V����(�k^ǔy��aЃz���4�{��l3�������I��{��I��9e��m�o��}�n�� ��{4�������5;뜗ƿ8_��XŻU�+|����_�ϯ����_�����b{N39���g�.�Cƺ��և�ٕC�|o���?��Y*�a�_�aWĴ��/��y���1���{��9C��<^����^e?T�dq?���H��#ߏT����rF�E���|�O��Vٓ�������i=�|��q!��6���POk�ۣ�kt��}AzX���:������w���
\���ezP�puOo%�9G#�`�_�W���nfp�@w�a�q+�I�Ͽ�a��N��>s����yN��h}��������m����tca�L�eq��]=����1�[Cvd���Y�x�T���|C�q"ǃ���G�Z����>�〼:�l:�W7�>�0鿯_���u��z�?�Ƨ�d~ �|��Cֻ��g9�?�������v2��Z��� ��<����e��Ȟ^�	�Ã�)�K;�'�x�7�����y�}+���9Y�����#ڃ/2]�g�׿��}O�����
��	��?#?�OfW�VZ��8�۱��2'鬤�<�J���?�S�7\��8���3����������;����u��LV�۶���
c,�;��L�?�y����O�<�Sفat�}����%���>��q(�{U�.�T}G���I��O9�n��3{_Վ��_�:^����U>W�e2�b?�-죫����|~��j�q�r>��?{����=1�$B��y7�Ϧ�g>��ˎǐ��y��)��r~�楲W�x��������؟��U/�<���=_�o��:�;}>�?{���$x�����)�]�՟�'�R��A�oư��:�}ӣz�#��c�_��]?j�*=����xԎ��༷}k��y��{h��t*������1��F������y���W9���Y�)�.V��������y�o��9)�}�ˁ���v(�ޏ�e�9���E�U�uZ�Y�����ہ�g���x��E~��Q�S@Q��<���ކ�b,��w�i������:`3��C��.踑O��h���7�"��{E*���l�Z�Dl��L�?<��cP����{��U{�ú���m�1�@g���}����p��ug�����v�Ƽ|���91�-G\��b��n��C?gvEuoI���{��������U�j��8��k��a���%p�/|7������U}>W���G=�̯�sV�z�3R�˿��I���9M8oy�'����U���g�ϳ}wŷ������:�B?Q��^o�a��C�����<�s��y4�+����c.�����ï48�.a��$�yь��%x����_���i�2��{fV���U^�Q�q�����0�V��v&�<�M휟�p??���!������E��P>�潊�,����'��s��E�g<B����k��w��+c��/ʽ{}�v��i8�yx[����o����%�3{M�}��OT�\�G�����۟�7���d��Y��íօ�[��|cYv�۔|�Up��x/"���)��3�_������v��-,g�j_?��j�����oY͗���3���L�_��K���b;6�i�䙇�w]�j'�bp��+��;}x�0�y���}����%�����t\��Y~����Xݻ��!\��3<S�}��q�7�g������#�1�>�P~C��-�~���g<�R�q��;e���ؾu��֟���`���1-~���\Q�����L��S摥�?��v�^�w������߸ߞ�U�������{����������������q��G�����H2ު݈�F�j6.?�R�q�	�=o�����ݳ��Z\O�����g�YpY����U�C�OoW���޺��:׾���>��򿷋=8x:D��c�8��=���S�u�<��ƕ?�f�5=?��|�^���S�gE�C��~����X^��?�~�6��l�C����}�ȷS�}zpV��Lu�]�W�6�j_V�+�sY����w������p:���w[��g�Cn.� �N��`|<�埇�g������'�^E�0^�t�3v��s2�4�N:#4t���0	�h�0�h� ��aPp@T�P@���zq��|��u����u�ʽW�����y�gW��=�_������^�V�Z��jժ��ʾ�~��p(��p�u��g�?�=<j��>�e��>�?�Wy~������ZT�+����U�gqZǍo��sZ�c��/%����0�:z��U��|fv!�[��!'�8���ؾr�;�5��xϾ;�Y+8��@�6�n՞�x����>��(]fxO�y����!f�z��u����	1o�2�;�_�q��e1~P������z��z%;/�tN�=���J��~��G�߯�g����~Q>W��/x���S���������؉Wd�G
<�{����p.�}"��+�&����i��P�}�O��7�g���)�G���qN���ȸ�罫ߒ����9n�u�^����O�y�Y��"�G���h}��%����uq��/�>h�[��_��a~�r����D��Z_��v��:�_��T~��/�6�~��l�7x^���IN��z|�}��n��P���������'�o�^d�x�_��@��U3���'�V������ھ���oI�S���{�M��9y���N�T�k������o���N�Z�SgZ}�1����طzm�����W&�<'r�m�}>����_n��!?�Wc�~�?c�o�-M��9�Z[�����rҚ~��3^z��ާ�v�����>ȸ���������8���c�R�x��p��o����M����)��/Z�M��֫x�¾k]����;��B��~�6����}���7�}��gyF�~����27.Q�g�ܯ���_�k�E��V_׏*����O���;=����������o��Ջ:ȝ�u:�y��~���7��>������<U|������6՞���]W��/j��'���B��8o=O[˜���s���Y|F���ko����a��]F�O��\��>a{s�O�����/�sn]���u�T�����x��|f�����'�st��U�&�i��p<��yJ�c�t�W<�;����5��_�ao�����Ų�C��./1��v���9
W<���'��3;�Wb�{�蜫7>)��p4���ۢ]�׼������j���i��N
S<�|�>�f��υ��	�u~lq��q]|]o��wɇ-���Q�!���g4?V��y��Y������;��=�?ÿ~IB���t�*�/s�ȁ��N�c�o.?��`�_�p�WU�7;r��B=��z_�2��S�U�u|����[ ������~Q����~�ҏ�;��Gc{�x��,���[�vſ_�GR����T��W�U<jN���Z�����F���J��=o�xe���!�O\.�,Y}��+[���?��M�o��x��¡���=Ü��~�����;��[�?�f}���Wh�R�
Їyuy��x�5�dv���-� >��Y����;�{v_
���D��}1���>�c��Â�/���	�s������a�4N[�A�o(��|Ϋ��!;7%�b߲�fv�����-���?�þ����J���?��O8﹢Κ�o��~\�=��Ӓ���Tyk֯��������K�W~�5?�j���[֭#T(g~?��խ�������?�?Cd�������f�[�L�+��
�<"�'=�vI�/cl7����2����-����O�փ1���������ߖ�n5�g��z��m�3pv�������)9d��m��/���K�}C��A�©��w�WS�k�£~��_@>�C��#�ʷJoTy�ap�9y��뫜ϩ�}k���P�4ぱq?��h3�q$�[�.~����[b�?�}J��I�����}��h�9jB��G��ϵ�/nh�uM���}�_�:��������cZ�N��`�������V_σ��ۊ'ÿ�n�#���P�����F ?�|<�Ә���3ݏ��5��^Fϑ�D�o��sđ�m�?{<goQ?
�g�g�o�#V�j��Ē��S�&��e���~���9ي����Ο�1�T����rS�����1��"?wP��N��3�̨��}��S��x��#M��]]��:e�O7W��M<���������[1�ׅ���8��l��Xk2��}����	���;.�u��B�??M�_�OrN���z���=�WY����!Ʒq{�����O��|��q0�\J�]���{�{�����q<1V�:_�.�3�ʜ{qY+�y��m@N��8�[�8�����Y�^7�n��!��o���y#���9�J��z 9p�?_�8�_��h<���=�I����L���}�_՟o48㜾����L�cе~/����|vy����g��횞7�Η�\=8iW����{Z��jV�,������~����.���^��1��}��K\�4Q�}ۍ��ūkV8��8b}��ٷŐ+�|��^��Y��=3����x5�������k$�l��{���~g{ľ�5>V��M\�X��H�g���	۩��V�ϰ�x�0�[o8�7̻R2���>9��,>�T/)�����bXo�t����CQ���U��/�ڮ�73����xX��
�w���3��y�9q�
�}|��S���>$.�w�=�G���8*���z���cq9���=UY���j����"?����8��:���U�븳�|@�����m?'�e?��g�)��d����`cyF�����a?��?9��::~��C����9osn�;���_��O�Ϟ���?{xV=�t>�?7�v�W��S���ܯ���=`��l���hm����	'ݜ��{�i
^��unu�*;tKgTtD;t�m^/��}6����;�.2�+���#�\"��qS�\�a^>7V���1�%=���C�ԇZ�[����Ǟ+�K�s�������ф�۰���y�b,��G���v~j�y������Z���K�$�^Ϲ����mg�_N���TmEf/"��^ō�>j��	}���^-������Z��\۪�f��/�q?����9��v���s�����Y�d�j����9Rw��}_r��)���������ғ��L�SnA��{�Y�*o��~3��n�N�R�g����%���x����#�xn6l�z}:/r��.ߵ�o�񷫸��b�%d���*W�y*�����U���]8xI�S�V�O<K�CeY��m� G�:�|O+���xt,+�+��g�񆤾�뭎��#����U���7��3�<�������XF��!ڇ�ȭ�w��|.�������{�o1��|x�G��qj��|���'���ot���m���R�#���1�պo��Kۥ>.�����5����}�S��*�W������5U܃�|�O2�s���V<�;���_Y��}u:�|
qy<\�K���Y���Q��v�3���u��Y�����;c��������w:/������.�U}��կ��M>l�jď~K[�mfV��B��v]o��?�n�9��u?"��n�1���⸧_'���׃>�f����W?R��A���:Yv��d��fp=��w��w����m���u�˹�k*F��]1Ļ��N�H������������ap��*������4y�y��	��7<>������v9^���8r5�1'�N�,�O�����g�������k��;����όU}B[�8� ���q������Wv�X+�}b�'���>�#g��_=�Y\��_�T�@D�7f~o�G���T��<�yQ�O�T�j�G�܂_o�x�Uԟ�/�j\����/�n��ʎp=:�������`qsl�6ޝ��K'�G��q�k��c�琶ܾC��{^�Mſ��W�hQ���a���!p_\�����a]�������V��?f�/kMc7�e��M��8����Ԡ?����8?_�p�u����/�~$�+xv�p�=`K�S��=������8��r��G�˺�P�/��i����.츱��$��=���9zD��b=Կ�38�O[�x����:G���S#�gv�������`��X~�_	�{8�=�Y<������Fv���ű3'�>���� _fȣ)��/������������W�zGE}��k���/r���C�@�}���rr�?���|���1~�
��OԼ&�O����}�����)��O�?j�O�r�����_�ut5.'����M?,`�s�z��W����L��zDK��]���Z����ju��v������̻�~������h^7
c�s������:��h�Y��گ�����䶵�I����v���#��|P}5�gU��#wأ�1���9���;k��?��\�<�����[�wA��}��S�ɉ�g���k��ј�W+<��<����#~I��-�G"�g����^o3���Xϼ���|�qΟn�����y�_����"V�k�0\n�#r������)����\�U3�u9���D�d�b6��ڰ�;��!z����� ��~��V��f ��EI}���\�+A�d����l���+tHǝtx�c�〞�3����v����Gl���oo�O�͏��y����j��/0>�T��@��C���kJ��-����������~�T����;�������򬰌Έ�����P��ٟ�3x�_�[��u?�g�g�7�}�����p?����y���秞Qx��������WmW�{{��~Wc��k��2��ɱ�����?��yE��ZO��B�"�Ͼx���4��}�r^�g����������&+~��~�'%x��T�bY7�
�?�����Y}�q�E���ק>w�������u.�;g��pI��/�ޕ1�',�>��L�9�ħ
��si���9~��g-�����E׿j������$��m��	���`ԉX/��պ���gU:O�<��Y�[�}"��]�ҷ��k_?�c������'�<����S������}���od�c.o���C�8'���9T��Ϋ-��r��R��G��w�_���0�wg�+���	��q���1��g��gFO�������dF}����<���7��II}__T�N�k��1��g�w��N��Vv�����վ*K�'@ޫ�	��W�g���έ;~�!�?ŷ
�Ғ���a��K���K�;���1�Gc�g�?��}����ʧ:]`*z~*���d{nߩ����<���ݛ���X2��O��8���Ku����鷸]��m*�W�9c�Y����~���׭�^B���}G�Sb����u���ݯ5��R����ta)�9d��"�N��<�jQ�c��k��o���{�+���y����_���w��dz�2��c��|jw�Zqi<�r��j-Y���*�6�~���
�s�����*ύe�>W2[���������O����Z���������̹�5Pýx��?��9�*��}���*���s	|��Ù�H}���o�	z9yl�}�:���m��W����W`��2��������3��~:���u�~�����k��u�U�����_w�g��X�>ws�Y첾�;�kן|o��'�sw��7k����W�O|w���\����+�S"��vٟ}1�+�8|��|�>�J��?�eJ�����3�3����ѣ�/���
T���T��U��]͋��q%�u̯��Y��e�}��a� =��X��G��Ѹ(�9�3�n�s7U������Z��ǝ�~��y��Ke$�k��T�/�8~<r}�e������ʄ~����뙻c�����oE?�pY�ƣ {��-�?�����7�6@�޻��z��1�OU8�|���י���/o]���λ^�^�c��,雒v�2�s���~����T��ՓN<��R��#����=��.X�ݭz_�����S��+9�op�ϡ���o�;���?��v=n����w�߱	䢤~�b���k��9bu��T���x�	�g_S���O�Oe�[�E,c�o�_����1o�kٟ�{H�N��:��{��P��g�����
<���C������Aݟ����kc����'�㋶�K=/���'Ǫ<�g�gM�!~�r*��Zo�;��d��U�T��>�)m��i��y��Z2�����e�ϋ�Fqd���R�i�^�a�m[?�q��#�*�.�U��ה�S��L�/�o���xX�:���Pɭ�Ge�2�)ۄ3O~w��O\��nȝ�[g<��3;���������F�����Z��wF�I�����W�,�x,��{�����{zܯZV�������~� �?��P*���r�z\���xBo�vY��S�?�ô��=�|�\��c����7�U~D������I��s��Ƈ�o7�7�v��"k��}b���6U�]��/�X�?�[���{*W�O�o1�G�#7�-1�k���/��ι�.}��걌�yO��}j���vF߿�	�����=5����h�키~Ĉ�xo5r�~�}f�U��x�^v���m=��V����	|yu�<�|v9?9�2���Y]���1�-;z~�N9/�rK���5b���}F�2�g�=N�s��.�<U}���~.��o�ռ,�{v���k�����1ȿ�#�?s�Tr��4�㮷����<1?�p�~��@<�ٱJ'i�v�(�O�*�ԛW�8��^&��+��P��?�p�����ϕ�L�3�z3
8����Ǐy�����u��r��V}W�?����:���;��Vx�x�U�����W5n }��nk���@�+����*���b��O:ֽ"�g��g �j��x��=�,ߪ�l�GA���_ښ�'�0�[R���(��w:��Q�x�����}p��k-�>(��I�����EO7x��7��mnܲ�7�WQ�iW<?M�x�{��I�VAO���q!�u�9���~]$��{�9w39�o��x���*�A�9{���cet�T���~~��}�LKV#�|��4�q|��7��zϏ�����|��5���g�߻i���W�G�;I��������;<N?ֲ���G>T�|����iq���r�U���)=|�@��_b����������gq:����q��>^���{�t]��P�<������v����?w<չ�
�N���*�?7����h��!Z�������'-��=������\?����K�;�����Y*=�|��*��f����q?�C�i�Q������d���ӊ��G&tz����=��|���0��L���ץ~n�����{b?y&���j��ww�-���y�����
���=s�ػ��:]�/p��Ϻ�pq���EJ��3�_�V�:O���`Y\��W��������5��Wzۻ>��&�/�������@�+2ΈO����Q��+��>��>뺘��8��rh�?�S9�/�k#G�[�̑�W3}xV��|�)�W�|k�������U?\iQ���}��O��k+�)�E����.��)\��[�f�,^_��v�_����	Y}p����9Js�s>�ׇ��X��E�����qa��M� ��aO5o���ᐴ��3T�X���t^�q<0v�ҳ�������� �/���i����n��~?w�~�f��\��2�����X�7��-�/cU>���+V����7%�W�ŪsU�_�������_�.~�xN��W�S��
����ߎ9�ݏǵ��}�Wr���s�y�����48�&p��E� ����σ;��bȷR}��y��5��0�>#�~��^���I����[�)\�=Ϣ���w�b~b����^������|9-U�N��p���D�3��+}=U���՞/ib�xtʱ����*��/����>�_������_����E:϶�V��R�_�ݭ�o��,p�s�����Wzs�C1��a�c�=�XC��0�z�Z�dz/�s�������O?�Ĳ�ڿ���x~��R�jG��:�
��er��ʲ�N.�T����ݯރ�����*��s^Q���ǩ��u��9�|xʕ���x]&W�9�08�R{Ȭs����+���sE�ƫ�������e�O��x��cW�l������w��%�#�����L#V��v���&x=�=����eF'��������D;�����"ω���
��Kl��Ƣ�?u���W~e������w��_ɿ�V������_!p}O���
��J/)|*������|a��֚?�E~A����������&p��ڝ�;^�}�.�i�c=���e�˝��T�S*?���g���7
���9�C���V_�v]V��T}����s�	���~ͣ��of��u���~�?�{��A?�[ןr}l�-��׫���9&s�1Uz��;l�8���:���������z͗��=�'�Zz��c]��ɓc�糸>����=T���8�:�S]#���~��y����o��Q#Y���^z�F�������s�ɩ��W�R�-�}h�|_Ggω��������f��Cٿ؃}����,,�}�{�焝z��1��7���0B���h�6�d~�������w�/��y���g
��n�i%t:�u���v����8^�~q��~�:H�[�U~5�c�������y�������7ڴv��qC����z�b��wƐ��s�oI��������T|`��R��
׸���̩�{���&n	�]�cl�X*9������k���U�~]��)�'�J��W���n%�O��X�fq3�?�i3���8��ɹ��g(����f�W��Gȋ�����3]~��0V�:�1e�(�yV�!ᴣ~����}�����<5�<��O�E�_�=���F��7#�9�E����:5���5�G��Y<�L:|�TΕo����_c����1g�	�=?�|Pz�a��븰�ͫ|Y��r���1���g���B�7�u�B����S�CW���&{�y����_���-Z��C���Y�/p���O��}�G ~�?���1^�3�z�pǳ�0'T�G�&��?���𺤿�?|Z��s>^�:b<���H��̡K껼U���֟�v�|�U������Z�u3ӷ���>����E�cޑ���i�'����b^�iw�r��S�ɠ���:.�"�+c���:�����7�'.��"
<ڦ«���3#?���uD�O�} ����jy���)���'Q�bN��q��M�-�:��q�3z���j��87���1����A�W������i�kz~����������%E��ī�H��o��v�^C,�8�3˘T���X��'�V��?Y�����cl�υ�A�W��s�	���MX*2�o���s�x���W���=�b�guߎ��s�~9��~=�üW�����!r����~d��91�_O��_n|P�Y���>eߝ��3����{�կ�����2�S������td�zs�����I������!�O����o�nJn�oT�ȝ3����7�.��j��[�#��r� �n��5F�}c5':�ψU~.�~�������|�`�"�}aﯞ������a�L�_�i���_&p�Q��<�2dh+��ҷ��~L��:O5_W��7���P����(kw��}h��׳�\�c
�/p��h���;�6�n��:v|%��
��j�7�.o(��L:<������ֿ�}~�ѩz���"V���N�ڝ*���X�<����B�0e�L�x^�=��^|[��2���8�7X�C���/k�~�;_�T��~�����BfO}��?�5���*>Wu�s��I�vN�yK���b�⯷
���;*',պ���,���h~��c�.���Q��}Y����G�~�����}"���8���R�^���{���o�0/nI�e�S������h\��'���z0�[�CTn�����M?��{��9�=?��g��q���_�W[����ض%���;b�w?c�z�����(�S��o����q��կ�z�cF�h^%��c���C�Z�~�u1�����ׅ��^şO2���8�.�"���^ޟ�[���x�	����}w���|�#��w���l$}�Կ���q�|��7dq~�A�c�����sѮ�ӈx�c�7]\/p���<����Q�O�<���Ǝ�2�/���ݺO������/ڬ����}��X�~�]~n��v�^,<����5e�l�7b��m��q����*�N����N?m/�����g�\�#y�����؏
|*^�x�_�K�ԟ���2�P�cy�����b,o���6����)~R�y��:Y�OV����0�� Vǫ�?�:Z헮���X�d��<v�ɋb|��z��ٽ��/�/
��?c��\u���	�Y�ߟG=W3?Ku�i����^��ٝ>�P���.?�l'�gv�(y>Wx�؞�kӒ���ݕ�D{��>�3<�/}���'�F>���>���=�����z_/�篣��R���þ��c�s1���/|xY���Ӳ�Z��5����� ����}U��3Y�ö����F>b7�'p͗��Z�:��_
g�2���>|M�_�.o���f�(+:y6i�<u����~���%������~����u�k�,c��]�j�3���߃x���eS����Sy>����'��ÿ����+����N��/cU`������a>�o����k�|�':q�9�e��E�t�xV=���u v�bG?��}RA�"�z��=��uzF�Š�p$���/�W<U~Kq.`�.�E�?g�z�<{�7N����r��ؾ?|{M�vd�}/
�\��V���+���?i?�}�J�����!�x?d�93�lv>�c�O���O�G���3uf6�欯i���Q8��z��8	���/2>S6������+?*������^��E��T5����g�+�g���I�_�!�x��g�?�r�9�1�{c�Vm7[G/��!s��9�|�ʯ��d��3巎�͗��	�W�TxX��-���1�v]�Uv\�O���c���I�����~��g4~�2�tV���l������Y���������9�g�j�o<���6����)�/cG��������S�������5����{������n���ߗ��K�����!{#_����z��cV����1���,�Ǚ���:G����X\o�} Y|��il�]�i%������{��>�g ;�;L:���ohG��z���콍U���5��sb���χc<���]|q�?�>?S��A���}W�Ը���:��Ď3�o.������*o�s~?�_%p�)S�^�o��<�{�*�	��J����_���}%��.W������W�gͷߐ��>���j���~����k�W���U�Wχ���Y��h�������7����������;gv�%�o���Z7��P�q�����,����"�;�����v.�Q����y1�+�#
��یa����8���䘗�}��y�&��v�>�����������_~�g��;���Xի�*�*g�Y$tj��y�����c<.�k=���R�U>)7&������YиG%'����{l��/N��v�U�����=�E���� W���? t">�����m���Կ9q�7
��e���L����L������dq� ށ��|=?E�.4z��5s��v:ԟ����y.c5'/�q���s���ܳ�~H�H�U�ۺ��Ԏ3�}���5�G�������)�����j��̇6�vn}\��~ �5d��3A�¡�/���.V����&�t�����6��j��|��кY����*�<����_b^�+"?���Z�{Y����R�e3r�d��ֹa��.+��N�;�ٺ�����p�O�?����w�c�_7'���m�o��Ö���8&p�u���������@�2>|Ro�h�����0�w��j9�G�-:�ԯ�~�ϐ�J�|�2n�������8���}Cϟ����;�'�=�����I��e��~V�V���2r{����3��Q�����_P��s+�|���o��V�Һ������`34�A����+|�{b�C,�X�{��9��\�_ʷ�>�C,������>�����=�냟�����X��τ��|ׇt8bo���d�lΟ+�w���="^����]�n��8=�����wm�ۭ����Sz����1�r$ 㐇/*����y^�]�y1��_'����Iߐ����|�1i��l3<�?��16��[����y��G���y��	���j=�~l�����������<�Q��T<,���ܟ�޺1��6��s���}�q�����~	x�y������;�;	J���ɮ��. �h��ٱ�f�Wi���9y,��Z/Tp���a�n�!��w�h������8��	�����R������f���P�T�����N���{9������Ύ<��}|F����u����^�"t��+�1g�����f��;]g�]޸>���_�T�F�G��{�3�(���V�ߣ��\�'�ܓ�9�|�����Z:ƅ�����6w�#r���k+��[�>�s�������@��O��9���>7���ysA�֧_q����׳j������s�W�����K�ݮ�T�N>^!ut~�`]x�����9?_�R(~�7`θ�Ƴ��k골|V��@΍U����ޟ���7D���R���9W�Q_28�G���>�>>�?e��q��E�������-�X����f���ߋ������H�/;|#��u�ԟ�.�棎��/�ϐ+�C��T���zo��q������f����ֿ��*�x�\�������׃�w�~a�WbxwݻcU�\�����ؤ_վ��C�]d�e�:��K������E1ϱ&�^���~F\������a�4�V�qU<�W��ø���}����Ɛ����/$x\r>��Ų0:I�2�<�j]N4�t|jg��܆�������?؁/>��Ml4�fC�͵���~��K;x�������i��\�/�6����7pF�UR�~{�u?�|���o�Ga�G���v������V�4�C�"��|�-�_�s�Tv<���t���7پ!x�q�{�Y��d�� �N�{I����Ie+�J}��/u=��W�߸n_O�B�f���=�L�g�{�_������E��g�O%��5E�����h?o:~�l�Izލ�w�Gp{D�[�����:����^�;M��3���}
�s>��ޫ�Wݣ�i����ո��GX�wټ�8�-���<3g�W~��g��J{���g����{a?������Aw����2C�����R���Ydz�s����s�����Z4��y9R���r@��y@�ĸh��
�̑�Ϲ�'{��jCp8������Ҹ�¹O�{U_#p�]�#O�<.|8�r[�/�炤>�J����/��ѹ�3���b�gأ��]?��vyϓÁ��_�ۅj}1�3��v�{-��wvG�~
�h7�< `<�pޯ���jտҼ�3o�ƷZ��;�?��R�ϰ���}#=��n������	=^��k���_���۱��V�_ǣ�s�~��s�
Ҝمlߟq�	=6³L������į����'�����E��b���j���
�c��Pk�uS�̧��i><��oS~��������	�����������2�T뿰���n��n�>(���A����;\wZ�'�����߻�g�����8�������k���s:�km�W�.��|N��tVz�p��E��[��Σ�'��xV��u���-U^h���M��G��g=>�<Vx��C;z���s�N��{�T��q�o�I��S?cީ}���2z��~,�rE�.Ϙw�v�5>����O�����}�!V�)Wy��§�g�l���^�>����42x�W�;�Sxe��?\5�/��p��ɾ?o���>��A�<��*|�_����sc��]�Q:��R{�q���~�{m��'��#1��>\�A�|q��t>(���������N9���>�I��TX�q�o��T��<w�K�+�bX�aw~R]<D�]f����&ŏ�=^��f��e�hÿxI�
�d��f���`<���}\v�g�<$u┼����QDnO���>*���~�ṭ=�D�����yb~�����3��~>��N���n��9}�M����o<��Zk��ˊ�z�
�+�9���������˺sY�.��K<�Q�[�׾g�)�g�,��N��a�U��6�����r�g����G;?���q~җ�|r����6���O�����/�����~�+1�~a����5Y�'���r�5�����������|+�Ϟ?05�2=��]��<:=�{����c'n�~��'G�Tq��b�7���0��ÑG�����v_�u~�t�>5��.����Uy����	��G�X���TN��a�g�ҷ�Bޜ����_�w60�꾥}�9��8��j��]V��
��N߉������N��U&W�<r���8\�'�̟���g<�O�_u�w��2X��+���I�>��8��k썱F��S�x�^�ϣŚ��?gx(����9j}��q0�ϋƫ�8?�����~��l�m����	�&-~]��z������K{}؄g&�}���Yވ��W�<���۵*_�4:��O��2����vm#�.�>�;OS���x�ng��V�:�4��N�?s�ž��ӌ��o�}<+r���.��w���^9�K�#��w���W��{kL������_��-��uG�=w�9z,���_ezk`=��y�u�%I}�D�'t���\��"���!e�����|e��.��Z���K�O��є�z]~��_͗���^��[�_�e7q��q'�Q����cE��^��x� ��~����V���9���������/Ί:)�G���([���3=�ql��d�}GѮ���+r~��ޫ����'���0|%��kN����T���7�!�
Ķ���OX���C�������[}��@��=+�8�[c�'��u:�ݥ�B���'
}�)������v�[��M�%.��׮�g����W�<�P�sgSt���</;��s�
�����K�eg6�������xߍ��	��WW����uAge7]N�g��<�O6z��ڮ�
�� ��c�K��;]��u�l �]�=w���r[��������Puޝl�r�r,ry�ΧT�s_��1�g�g�?7��j���mߟ�u��y��O����*���p����Q�踜��>;��5�!��9��P������<�5�q��z�c����[�xCcʄ79���p�R�a�?sσT���s��!	��a����I��<Z��������g���կ�N���ũ|߁�%=��׿��}qAO���s:�q��?C�b,��9מz����p=ϥ�����ö�����q_����U�������@��_G<����;�'������>������=���(�Y^�y�9�������X]_����l��F�݈�<���4^A<�;���mV�H��p΀�������+9����G�����N�_��O`���wW������Wq�*��׹��p�@����q����VE��E�K�x/���S� ��[��������Lg��Ͻ��.�W���Y��i?��֯���_��p�I��sc��o���D��-�S߃1�3,���3���OξM����}�e��ؔ��N�֩q��������Cu���%���v�-Ƣ�$������k~ű�xW&�o�o�O�W�\=&�s��G>?��ܸ��<��9�}z��f�S�bw�X^��«u���gށ:��wE������=��xo��;��A�oA�d�;b|X�~W����c1��4�|��?��T~��F�������O�s�|��c�i�`]�yK�S�?�x���9��R��9pN98xo�ƙYo���<��۪hZeO��\�\���������%�ݟ�o�$��z��G��q0�~��y�l��ӯ�#P>ɓ��d��qaq����V�o�虫�]WN�_ő�U��+=���=����*[��˲?�kt��s~�?c�~X��:�P��C��.��gN���*��}�>���~,��G��Tr�|n8����OQ�U�U�S�2����3N���D��Y���X�m�o�7�?�L��P�����~O�"V�}|��hl��o<]��ϭ�-1^_����[����1���y��%|����?��g�k|�WߏI}�"��yq����7�u�AiW�����7�\���o	��[���bx�|��l�����ɑϗ�U�* ^��e��p�w{�=rZ*{��kY�������5'?h�r��S�?V�;�Тq��츿�}�_��^���*����μЩy>��p؁M�S?_o�zX��?��MѾ�oz�X����ߟ?���5��?��R�'z��c�7�y����O��a�u+=����k��l��*z.F�bǗ���e�Q?�V��F_?v��_��Q�e�*�+~�GY�;
��lV����Squ_���i���~X��N9�_Z��i��{�����
8t?���؎}��n�����/�hV숿��S:�<kr���/�g~Cz�1~/�f�s4�w?O����[ǋ�t9�sA��>������<���1�3jO�����M�N$�}^�����Tl���w���/&�����?��~�����kB?�؟���yT��F�
�������Gc��z����);_�����[P�m1�% �c�{
*;���dv�m~�}��m�/�,{?,�s}���~q��>�gF����?��a��Iu~��¦��hz��G74���M��.Bfo�<>_�So�]�9����e�����z�@���u�_]�)��@.D/~�}l���m]��]���\�<���r~ߎ�}*o\�c�����y��gD�o\�K�x�;�0%����ɿiU?�5{MBi"�ٳ�-��g|)��}(����:D���������'�}�ϒ�	�y���/�y���
8�:9 ��(�?����$���_���)�z��UV�*_��b�>Y��o[1>�=e/������^p�P��9�5C&�~�q��y"w{_���Ϸ�ϖ�O��1��]�޳�6�Nx�qE^�Q����:;���V��6+��K>{��q�����C.t�e�Q�C������O��!+}U��3
��?#��U���<�����z�Z�Ew:i��~����7�@�����u��+�3�}6cU���08��b��T�x8=Ϗ��wKR?�Q�܏2���{�M7T��� ����s�}n��|����Ǟ�g������w\g�������!��4_i���q�`�����޽��r���v=~β�os����{ފ<���j����ӣ�Wzf7���ݏ��?о�ZS��8��_���������*Óѣ��L�[l���|׸�����C`a�j׾���u��{�0/^%�c1��X������s��_�X����-�Zb�_ݴ��_׹zo���ψU�����S�~e�(7��\��N��n��n��������s޳|�}7U��CΜ�9�e�q���|c���]��׻���7S�)?��k<Y�Ѽ��ߧF��qT=�d{���MV����e��/=�@���ó~U�����g�&��Ι/:��>�ӣ����tz���c�Y�}=��ߩ>DY��>d�����Op�_ӟ��X�̫89r���Iԃ���OM�<�p�� ��3�w���8k~ �{[�<[&�+�����=���X��e������s�9ȯN�B����ݜ�@y���[���5���M��{cX7X�h����k��a�C��h�������L�׺��j}���h������s��,�U�7[nE�g���ӯ�	g�Vp翶��+=�eƺ~��x���1η��{��̉+nŎ�S����8��{<2�9���zL�r{8˔��%p���S�1��,��E^*�Xތ1�O�����~͏_�瀏|�������_e|���"j;��7��������v��{��z�e��y��{Cc��g|���*�U��sۭ䰪q����1�<���z('�Ū�̳zսٙ�'���ʡ�'Rb]����W� ;���<�e�� �̾8��Ϥ.�s�8����>T��{[�xiL�]��w�7�[���ܾ��D�j���p]s���Ocs鏘��_�a�y������$��o�?�>����_���9�����Y�y����/p��T�&�������|����G,j3�S���g�-�W@8��E{�-�z}�t_��i��q�1x�/���r(���~�}��B_��S��y���p��ˎ炤���ny�����W�F��q�X������^�<*�,���*OX��9�0��;~/7�}���6A�'�j+y�W��B���_>��*ދ���;��U��_���2[�峭;׬���V����x��~s�����I��~g�+_���>v_M����ռ��M�sZ>����ߛz.��,��=i�]�n��wB���7F~�#�����������9�j~�v���X��2�~�1��]?@��z�4f�n(�����#���c�J�V_��w�mF����O-��>�!��[ga����$�ɫ��,n�|�w�ߊ�;�_�ϥ]8������~N�"��8��/2}Uō=�R�sQ<Y�����n�yn�E�����'�w�O���{�/�|\���Ϩ�q�呪lM�|���;&���E�y}�!^��t�M����n��N��u�7����i/��g������A�.���뱸"V�5��1�ߘ���Vd�í��!'�&�F��~���J��8�^�9���ݣ�B8}-���Ga�`�dt�D��:���U�N�9W�<y�<��95_�pޭ�WV�R��<��CϫV���A��Lh�_T�Y�.���)@��'�s�̉����NϜ��
>�t}>'���E�Wuߋ�w���<h|�v��0ծҗկ�w֝�����Gx������z���q�7��+?�N�/�����닩{3�y��S�W��>g�]ᐙ3��_��y�Ͻ.���\����
�O� ��c��%|�|T:ՎT�$��KY�,>^�z]ī_���~Q�2��GT>_�ׂx��������C�5��ڧ�i�K���ǂ���_�y
����p�P~�h��|�ԧ_�ݯ�g�l���n5�R�/�uS%n�4��3{��W���N�ݯ�*������펇~���Q�u�:}���Y>��@�	x�/E�����hc������Ӥ>b��wl����+z��0ʜ�,��������=�vR��>9�|�q<M�_�zX���U�K=wy�����/�Y���u[�i��]�W��3b\������u��ˁ���=�8�x���y��b������<��+�:��{�o���w�����[��^��(�z���@�?3�y������!��G��\���v��{��7�z�!��o��}�_�����[|s�����Y��7�)�UN��OC�|Sp(�*�T�T�0��=���#:�M�uC������ǋb<����z�|����:��9�8f~x����N���7~� ��7�[�*oW'�d�A�9���	G���)���v����k:�:���ӥ�z����>��X������O������9��Ҏ,c���QȩzU��ï�w���������+�CP���=<���y��$�W��U\Z���� �_ߛ���#���?̶��$='t�߮o�>���O�?Pгn=��9���;�x�u��$��<���O������X��CҞ��h�n5�Ό�8�ڗ������b\t\�;�w[����� C]4�'T���՞f�U:9V��:;��A�s���u���p>/�yW�!�;������U#V�`�2��Ҋ�ԕ����2=��EUө�_��^C�z]ţy�����=��a~ x�~�����w��5��C	�*~V���.c�<x�Ϡ�9�='��p��*������0Ė^,p�Gb��y��=�������Ϋ�þ�O��w=�7�0�տe��L�����s�/��6�g�s]����`��K;n��ˤ~�?��yk��[1���<�����>�|`����sߏ���k*������G��v<��h߯1<J�«�n��M�?W~C��uZ�W�6����S��*޾Y��Ǫj�Z�Vx*8�)rjOz\R��Q}��y_K��~Ե9W}uI�c���P�jowz����
��[@ސ��}�:�,�wy^��i3y���J�����S�<�a�~��{����'zs֯*��Ԃι��uAfO�{�\�O�/�������n��89|*�]�G�������7�����'��?.p��A����+b�>%�[���;����ƣa����_��祝�i��r"���^�i��d�1}_����a!ϧ�����8ns��wN<J�*�?<���R���؉�}��on`����l#�,.��<u~p~����5x�GaY}�����Ǧ������M�1��X|]�yV{���|g�ϕk����!/�,��IY�*�iK2���p~��vG����tZ��g�^ ��k:�3���y�~h�]5��I0�/�H����њ�����Ʀ�\�2�5w}A���鹿���q������L�Bwf��u��*���k#��u��s���{��kh_�}o�p�o�q]_���v�﹝��U�\S�Y�;�4?��n����/����fF��?&��OV�-���5��K��ٽ.l�?��=��'�>^<�z��I�_�%��� ��P�����N�f�z�y+�s���um%?Y��\��t:�������W����S����9�xc��?;����C�}W�ƯK}�O;���9e�����9�/��T����W���*P~η�,n�/�ϰ���Q���|i�o5�l����q��9oQ2y��6�m��N�p��;�7^���1V��v�|���{J+�N�+��TI���|��c엪����_��������{E.W�3���y�O�/?C�+=O���J�@��{�k��������3��M��}�չ����~~��G���������ya���nGX\ N�sן"�S��گ,~V�F�0���'?���8$KW�w��ǚ?��}�n��9�띪�'Qz�}�:���׃�OA��g��si��}=��1�z�c��It��o�>B�A?b���sV��V�ED��\w���+�>��7�����>t��s��{Z��k����0�G#��>�V��V�=���m��k?��/H�Y��O΍�=�g$����������j�U��}38�"�e���/�?��D/�����s}��$pow���Σ*������R�3 w�#v�y���!������������=��ú�a	�p�"���)�,gyA���������ҏ�=�>5.�x�g�qW=�R񳺧��j�:^��~4l�wE>�jG 3[1����w~6?y�}�̆��p��� ����S|�~���e!�m1���7|^���Y��͍kA�������]}݁;!�����4{�ܾ�u�4�4���}JBu�����w}��[�֩���_���9���g��9=�����m�7��k�������c��W����7q��9�;cM}�[�����V��G��j���G"?���n�>��$?��k\1���׭G28�&\�������?��z��I�u﹈^���,o�����2=rN��狤���y�w	�k;M�{Ì~��(�o��A�������<%���+��}z�X��������$�c1�W��}�o���
=O������cQ��<Wv���ʧD}O�����5I���P�=�8�'�?�y�P�����\���_��T��s:�<����'ۿ�8��_u��?���~���F�*�������˴'[}�q�z|������z�b<N��~U�����3����24��k:n��+�:�|�L�(�ǎ�+t�E����`p����ܓJϯ���s��Ã�� ��EI�,S��`�O��~k���q���;պ��l
~�G���ª�u\w���Ѣ�W���F�Y���*y��<,m*�9�2�y5;�=�o���t�A��ˍ�=�zl?cx$�/��o||��s��}�����0��}�9�8���ض!���7��ͯ;�%��<s��+��G�.����Ç&x�o�<�|*��qq9��)����k��������3�vV�P���6V����6��,/(�����ߧ�Y��>�U�L�䡊�N�q�X�+���o�<�+�;=���������zf�.sX����<7zK���O��G�=�����u�9�c�b��/�����^/�/����~�_Z�����0�?+�o�t�|}��,�6�x���.�������
g�����\���������l]V��ݮU�;*<�7��e�%�}����q�S�[�� D>��ïu�0��"�|{M��?|T���g�3o����~"�9�T~ױ��D��%���~�n����u�����>���n��Ϛ�ߟyަ�\��������2���=w�۽��8��2%W,����lS�����;ɛZ4?r��46��}��(��m/�`����GΠ��s�♐Y�o:��=�����%�Q��G��O�ǖ�������cq�G��K���r_;�_���H�V���ռs��~.c<_���w�_v�#:,����93�kz��s��ޯ[<���՟���3;-h�C����,-U����ў:����n��W���)�~��?���q9h��G�O�	���S���b�Nw����������f��w���R�q ?/ɲ[y���n�4�J��7<��+���!��AnoMc���k��R�����_Ͽh| ����GXv���~!w�$�w"b����=��[vN|n܌�,�S���)K�7�\�yU��x�'������{�N��t���?aq���a�O�|��������\G���c?g��پ�t�}.��Af/|}M��qj��~����yh��6ɻX<����z�OY<%��ƺ}��Eϩփ~�IK�'�����x�>�>�ݹz��w�O��_�/S��>����!����]�q:1�.���g��Т��|-���8����Y�<�����<����!�sϹkBV��o�Ϗ��������s�Q&�{�ϣ�.[�#��4/8��Dm�3��1r��c��~�PǑ�Z���Po���}"ů�yo�~i9!�����z�8��/���,s卸���]�Eu�ҳ���zpǯ�������q�o�������w�p�Z�|c�ܼS�e��Sg��@/깡e����"��_}r����s_����j�x�Tq���X>�a�Y����ѯ~���}�N�m	�s�p�*^����y^���jwN�W�_�aUz#���z��<7�X�U�����;��Yg_�8����q�D�����|��7�n����bX۠�%xܟ��;��/��W4N��n*�����n-*W����u��}�?#�Q��1Ńx"ld�Ǔ��-��÷bl7+9��H�=z\���z)Ã�E^f���y��f�G�4����~���y����tޑЩ�����SrUٝ����M���=.��v��[�y�W����bl�q��b�qd���G������g�ks�y��7Ī\�����8\��|���,~�N�-s�,N'��=��Q vb~�C��"��4�~1��y^�����2_�M1����6�:�U�1�~׽M��۹3v��x�����?�xhG_��Թ9�O�A�7��M�����m���B!����Z'�<@���
ȗ�K��ޡ����N��������g3F�����D���4j�����>�H8��]�g-��a����<W�q'�WP�|��g��=�7g��@��'�3g��p�1ǟ\��wF~?���󍼻cXK}��^֟��W嫨~�:�8�{�*���38�������g�U?�%��>O6�����s��9�:�����T�x�9�h7��ϗC�_�L���V�s^���C>��5z�߈��c	�nǧ�E.blO�f����q�|���3d_�(�oߛ�q�W~���q?��_��s�J\���k\��gfr�~������=�h�.��5�Î�;�n�=��6�浾?B��K���1�
<��Y���*p��?;����?��B���]��j~�ް��_�OΑ)9��Ϯ��?c�q��g{c�{s�S��(���K�~�Y���{�`w��8�zG���Wy���8��wl�~���.��O��b��s�ֻ.����y��y����7�'>���|J��/|Z�o�ޑ����t=�B�3����d�+~ʖ×}݅��H��t��;�U�p�zz���4_E�/p�q��k��,�������I��{�ط��R�/���{�����-�yr�{���	���?7�˲Y�΋�a�����{�\���_�	Yo�aS�N�g����:#���!�4Qh:l��1~�+�����{�*>�<�OD}K��<���Ot]��+�y.:�}Fz�dF?��#Q�p�ε4ሏa=���S?�G �1��Lo�~㹂��_�|j~W$������Ό��_�O���O�q��?�M� �1<O�����}f�~�$��}s�����tV�?��Y����U��C?�g�����mW��{�������R�~����gƁ=I�ϡ�4�'r���\Ɯu�����_ŝ6z"���ϵh����~%W����	w����yB�z�ޜCVs�c��zN�ZG<C��8�3�Ų���:T�C>����4���N:O6:1/s=��V_��3�_�5��w��?ip�T�+>(-
�[�����O��+z�������N���#�͟��r;[�W��g��jw�<_4�<�6�i �D�}K�n�\���W��z��w��|�*���p�o(���wk{^��/Uϋ?V�ؔ~�yqM��d�ϱS���E��?_��/���N���WT��錢��Q�>ou�o���q�������R{�����x֯j|]>���țP����I��6�!f��E��|T��G�������G���hA��{4U�a��_�0V�w�=���������^��f��~�ս/����>��3V���b���^�{�6c�g�;�~�m������x��+��y�Y<!�{�oW��5�/�gGc�O}EǁqyE�gݼS������=���=OMyݲvI�f�g�����Q��Ǯs���v�Z_{n�/��?<�A8�{�f�נq!��^���}r;U��e��N�.��X��W�/��NӍ1�ר��5b6z�?���A��`/�6v'W�}����=�_�?��)z.����n�Q���~G~b����s��N�Q���j�Ry~���=ۃ;&��rC�	�|8�^�y^�ιߣ�`g�3b<^���@v��g_��;w�{Y���Ο�F�<W���	���G�����}O�����64�=�����L?��y�c���f�^�g�{u�����Y��s��n��������8�2]9���n�I+�������-U�Z'��1>�������,c����M�7��E�T���U�7�g8�?����z��U<_����'���t�k�y��O��7��6�����鿪���R�[�do�����o�-��Y�鯎��~������|��8�/U����/0:+z*�������G}?؜}@�G�|���>�����Ѽn�O������>bf��xQ���~
�7���}[��11o�d�Y�(�Wvt۹I�J/q�2~Ή'��}���~�}�o���_|���V�D���q��I1�4���B���o���4[�}�E[�Y&xx�˔���$��P�0���;��o���]8;u,��j��O����:S�����iZ
��t����;�w�p��[z����=MSyqߠ�z���q�ۜ��.�gDNF�/ex|���Ӂ�W�H����7�Q������3���Ks?�:�1���}�lsn|��9��?ם�oB�2����xBv�������lȞ�o?��o+������W�\���sjG0���6=?Vy�����!Ng��������R���<��a��"��u�����K�(7�v�C�RH�M���}�su�0��oI�K������̉�n�����w��>�����t���q�1Λ�?O}�|�~��Mݷ�_���l�7�����^��|r�_֚|Q#���O�9��kU����T~N��w-����������6>�?�=��9�W�!���iu���j�����9��{5�y���?D��/�-��{,����Ezxw?�<_}#��l�?��6�뼸�ׇ��}��]��;��<Q:�o_w>�Pg�fp�:1��!p�e��<���w/=�sy�⥄�>�/N�4�՚�S�7��������z�D�_J�������v�<����1�5�u��?��<����+����r+��'O�ug���޿���;���9���N�O���ɂm�e���<h����2��8R_��x(�� >���0��ׇ�|ć9�u�w)�_F�~���+̣���.��/�����N�לϚ'��aҩ�YN�v�����o������_��}���S���޷�c|?�Y���}"��}vys���x��?�+��f^������k�`�y󺂞��_���{��pA��^*��j�ل�67��/8����_��#�w��g��~���3ւ��m�w�<2��:�y�<��3JO��\Å���~춬;F�OTz�*^CO~e*��2�]�W
W�����!=�nw?�:W���u����m���/���\�����z���o
\�;s���w���O`^�2��R<l�^���7��L�ه�_~�gt�o���T�g|��k�_z�YE�ؑ�5�������Ū�ΝSz�҇���ϧn�jW�X�����{���g.�0���X�3��˄N���wq,�����[����P(��).�������xY��J\s�~Ӝ|!G���<�W���Sվ3�}��M�{
����:�5t���#�<n��n��5�J?�@x��א�rCBO���X�����p6��_�u���Zg��]�wn�� ��_�H��gbU>��J�,�3��<%��7�a�uʇcx���jÏ��r���{��}k�Ϲ��_w���u_R�w�L<�yI���z=�Wɗ{�;�践�~+⫏K}��\����ߪ8p����y���뵌���~���w��1�,�]]OQo��e>�����?��,{b�g���1�yB��x\Ǎq��C���磟���6w�3:��5�yaƏ�L睎bh�G�3�<��~���?���c��'1�\-�g�|�&�%��E����*>P�ɹ�,�7��q���FBOeǑ���}�[�~ǙI�J��Vԯ�Q����ew�z*��^A��s�h�0���<�X=w����sc���\ũ��|g��@����w�Iyu������ϙ�^V=��#�_����%�?'�e�� �Q�����2��yvO}��u�d�:�g�0z���^���|�|�}z�'?m4X�F����Wy}���sU��ý�w�x��W{=؅/8qy^�꽯+ڭ�S(��}Y�{�
���'l��y1�wb��`���uz��KL:*;��syW�x�k���K��1O���Q_�S2}�����hk���{��%�ٶ��F��vm]�xT�����޼�����r���R{��~w��ۂ��	��o�z��;(�~��A�S��L�U���p�Г٩�v�۞��u���~��ѱ!s�t�gD.�:.ȫ����������*0iw�՟�#Տ弮��<ؗv��N9��;��P?�'�1���cx?��cx_�\������p�3d�_F�殃�/�N��q�Ÿ<?�S���O��g�{��qo�?�;�lJ�f�V�}�����_s���3�{�8��q��޶ʾ8�U���視D�.s]�W�����,���~�ٽ��|��!�E�ݧ聞�]l~/4�Q����^��~h�3m#��c�G_��^��O�a�W�/�8�~ko_��������T�Q�T�o(���C�c�qsl�jW�9���gv�u掯�m���<�,���9؟��?���~髶�S1������]���3��}�ӹE��u=��}}qG�=�{�ѣ���{�_b�W�������m��p�7Fl5�:�����a�f�X��JOV���Wu<���'E����B�>e���d�e��ۛ�F��fe��|�zG�݅	��kQ8����J���b�#�*�J��G���_�᮷w	����sS?G�<�a�a�o��a���|������sVY�d=���,#׷,�v.���1.�W�3�k�T�]�?u_����}��g����݈\o`� ����k��d8��W�v��=�?��z�D��W��ty�s
�w��U)���<�:s+��!ߪq�xK��	�o�0������.pg�������{�;b$��}N�onl���:�7��^�!1�|����Ο*o��Z/{�H�OQ��V����~�A�r����,��1�+�{���}O>ߩ�}"��p�[������s�;����Z�78�\�ڗg��Z��&���8��sc��,�*V� {���l��~Mu>]�v�ę�ߝQ���~��)�����|=��~u~��I�K�J������ϳW��,�x��_8</c�sI����]�S��������X̾/�l�y�}���}�����_�U�D�k�W�����"��'��;��ů*9w{���AWi�_׭�Gׄ�����FO�J�	Y<.p�����6����X����>+�y,U�ا�\�EV�;Z�����M���x�����U��y�'�N��#�������烷����/�6?�a�y�\�za��Y~7�o��O��)z��S<���}�l>.:��P���ĘhR�������/]��>�]8�����)�j�]�U�o�W�F�3F��T�6
<��3��3:�_�W~?�_��ύ��=ŧ���O��=*�<��e��o��R�[���S����������~8�y}zOfw���,nO�����I��'��3���#�,�ݟ|D�_���滞U�������@�/r���q�z�޾��Ñ��Y����;��[%W������O����������1��E���Xȯ-���<-�s��2 �����K���y�Z��
��l�e��(�ߪ<:������+�xHp����X�P?C���>V��������:@���n�qv�Wb����h�ʡ��=7��V�}���Qω��R<o�ង��=���R��z�ڏ����}�+=�J� ~������X�$���%��R�|j�f�cQ�kP_�w]"v�|����t���m��O�E��ع��I�����ո�<sܗ1��,�}���G�ǋ�يU9g��{���Y��鿣?#pL��?�)ׇ=>�#�B�$�~�jG�m�q������6��ƥ����__�_(�sc����+�:���~*�z���U1_�A��?�ޕW��;|K������k��x_ct���j?�hk�GǪ"���_��3��Gtxu�ŇuvS�c?�m1�|���?~��:�c���� ^���v;��s��{J����Q��}�9y]��������.l�O��ت|f���슟>��]v�Tu~�����e���c,����~��´(�/�0�qݯGNx�x�MI�OE�O�pF���W���w�@� ��g
|��������wU���|0V�8�wH����mD�o�]�@��5�������s_K/=�ԿX~7%����Hl�#/t��.���6IGfG"V�w��}�F����o�z�b|���ӿ�s"*��.�\��y�*���z���7�m:����y�~г?4.�[����N=�����w�Q��>����ۃz\W��]�u}��n-�#���׾���o�W~!V���6��W�4�%"�������'��GG;迃	~�-��\Oi���ol_�D��ԔX͗�}^�y�o1>@�:���K�н�?������k\]�>�������pD�k��r�ɕ���l���F�U|��/b<f�g򾫹�Gߗ�^��X���_�X���9��������oe����:���7}w���V�N�g��w<���Z|*[��y>ȣ:\���ƶ>\@�v���U���ԼJ�����q��[�_����x���ǘ��U\b��u޽:����_�Ag�w�|���g�?����>^����c�#Ɖ�'�������ĸ�/� �<+���h<?���:4˷���xޚA�n�䣟���x>6���{6�~�/�ā���`���*!�)~�5�o��d���GG<����o.ƯH�JO�{c5�P�����������2�Ѝ�O��;�I����I����zˡ^�(��Ϳ?��Ž�\���O��~�яrI��C��.|]��8Ce����~����y������o���Y�	�_�]�{�NN��>�����A?kr�������#XFO�Z�g�Ϝsmٺ�����Vじ�wA��p����R�ŕ���1X|OC��R�~����OwC ��X�l�J}q���1��G��_<�����;y,�[�ϭ�X�����z�z�Ǘ���cU����+��?Ҿ�֛�7pf�k .�I���ϑ��~�A�y�s=�/K��B8��e{���+������a����۱�_4<�o� �M��u�>�������}m0���a'�XO�d�����{���p���=?y�ޣ�}]�	|���ݙ�����ѣ糖<ۤq�'����Ѹ,^>�����c��i������y[Wj�C�1u\*{D�q��\��+?���mv{�^KfX����!.��P����˖3�aq�1?���]�qx��B���C��������qa?}�\�-�oO�go��W��l=�r����ǁ��x,|��w�~c}~�Z�h��]R�����<���v��]����9~��Nm|��}e��=�ٟ�'�l���3:����]���s�@��z~��_�u��<����f�_���ٗ���_�~_o�	���tx�!sR��\��Zt\\K;�!�W'����vu_@ߗ���@���_�kc�����"V�{zS������Ob����9,�_ϫT����:���]�/�,���V�qy`�����4�����ΣU����?�r=�^�����qWR�����g�j^4�n_�g�?�?����;�Xi^.�^b�_����]��?r9Q�$����1�gnl$(�����jWq<��e��ʓ���yz�?������8�{�{%��������k��'�ڐ5]G��<�GI�n-�����1_�Z��^��>׺�Y���S�J�������ޯ*�T�Sn\���s)�z?��)�XG�]��=?��֕�M�q9�߫}9(p���yb��$�dOӏ'�uˢ�v'��N�K��z����>��s���ՏU�Z�#��s�Gc�_����{-�ϗ̨���n��i_��'�y�{w����g����� ��A����g�������c�W��ҩ|f�s�m���d?�W�'|L��p���|�c:~]w��Ô������RW�̷�q�|�,����{��8������R�Q�~��b|/�6�=��^���j"������SϏ��翁?�C>3�8R�Ǽ]��Ǒ|�u�}#�G��5�4۷r?D�.?��O����K�
Կ�����p�)��@~�s�v��$��S�z���3����d���;ߑ�'>^������a�wS}xr�;�h�������Sx6.�#���D�%�_�9�^L�q����s�˹>aqy��kTo�ރ������>8牟�־*������U�,p�a��x���d�_]����w����~i}�g=�pS����Tܘu���s���ɇz}��)���5�y��r?��%�7�]��j/��܆����T�1k���{,|�0�C%��?z��I��|��m�����E��8�1�3���N��5�7���,~-��`��+=_�O�~��7���`���y��>����O�����+�v��&�FU���������Y�:��(�7��ώ��p�Zk��o�ꇳ_�k��c��-1�?d��a�zzj�O=�����Y�z[0V:.��C}�����wA_���c1��k����u����$m<�ǫ�
qv�#1�q������������� `��uӅ1>�	���$|���*��}@��ߋ�s=�9�rnz{\@ˉ���{$Ooa�y]�U�sk��:F���4�/�'ߩ<���!������t��b<�,s�tG����"�5}M�#����N3���+�����]�:�^_�J'ϩ^��,�=%Fzl;O�1���|�۵e�����x�~��?�a�8t|����ޝ�?�}4�Sr��ͷ+��}��:��8���<�mvn�>�ʳ���E���������>::u�����ǋ����a]�f���{��z��������_kQ8����0ʃ9�����������m�<�9���N[���|V���u��9q�*��m1���$���W�5.7G�O�������m&'���^Tq<�/\^�?o18�1qNS��O��J����k��O��~�=0!����d|�����3��-6w��7Y|�����=���������@�gn<~0lWӣ���=���c��5��'T�tX���"�׬z_yu.{*���Q��ϳL�1��� i�������ƓU���K�=6
?��%���:/ԟ�>�2<�w�7��{oo�^6������N�WϷ������}���������=�����CW�vaJ�$'��~^���Ū�U�&N�C���1��?��G7��;uV����aq�뺻�G��}N'ֱ��`'�-���s��N�b�������7�*:^�S8�e�u���y[���|~���ܸ�9��U�������hN����?�虻W�k1Onn~��A���?�/��D���X���.���������������I�\Ϝ-���*1��ث�p�����^�=YC���3���dz#�_��]��V�!�{��1��J��u�5g��d���p���+���b�>�ކ^kszqs���W�D�Ƿ�(��u}��1^��ul��9P࿪�C�ݕ=�1��Z���eF�Ծ���|���q�w�X�`ˏ�X�(ǯkNՇ�ȳ��@��Ԃ�u�����d��ft��_�;���
^��M8��uyDY^����Z������4ί��
�Q���7��{�0�Gc��>!�C����>kw���ꇓ������M����_ƻ��N����"V��������ɝF�Gו���`ow3\fx��׃\���sm7g��R����'p���<���Sz�g���鎿�|���v,m#[G�d�B�G�*����3'�}�~����]������u��#��s���!��g�;�kv��X�����o�u4��\�G�{q�I�؏�s�����t��c|�+S��8�=����M䧺���c�S��p~���#��ि�Ū}�zj3i7b��@Ξ��<Tv�������ύ�lC����Fϛ:��/N����������ۮ��9[���f�1o�����}a/�a�i+��pS����Y�=��?��/c5�D�e�u��<Hĭ��{cgO������Ӹ�"V��[W��\����&=�^���P�0/��?�0�}<��qx�����Q����/�:no���}��ԇώ�bio,�	�ǥ�l��!�5��`R��L5�X�]��:���s�t�ev$���=��D��'}��7$�Q2��k����*�_��}�R�7R_����*>��OX�?��夺�I�Y���?��EI}����O����~��y����[|nR���S����@�͉_����?�߲�;Ǫ�a�m#�u1���gQ�+<�������=/�E�|�>�W�fv������X�#���@�4��gX��1�-���J��3��j8��˔~��XQ���C^&���'vܘ��ڑ9���+�{w�� w�DQ_���qĘT��+ݷ��������<"�v��-cX�͑g�3�3>T�=��g�e��j��N�c,��:���ݭ�&�V[	~�3밇�X�U������q���ꓦ�.+\�iQ<��9�/�_�������n��c��|���}����}OoJ�D��^�s�G��ŧ�5�����۩ֹ��WTr��q�z�A�-_�뽢�D��-��������w'�}a�B~w�tz�}p�y�^۟o������O������������2�<��3^�/�[��|�9�<��>�������Q�����C�ԯֹQ�Q�z��U�����ڊJ�����q8'r�i��N���V���o?-������_��/18���O������vgq�,���p9�>���6�7�s~��;�Z_8?�Ι���#��8���^��cl��h��
����4_cqcc��KE��;c�O��X���~U~��e����q3�?���o=W���?�����y����C�?��|�u�\���v�������R��
���U���o|j��e)��}X����?9��9��8��>��]���ev�z�������7?-�U���:��gw��K�~�q�Y����G�oU��bx?�gt���^���׬ѫ�C1̋��ۥ�{T"�Oy�xr%Ϝs=ߊ��׾:����-�v�O^�A�?~�m��O��e1�s��]��+c<�="��7���z}�v«�
�����l��U�����c75�[�w�[b<.�c��*mW���>/�7ͣ��:蟳<��e���,����JJ�i�qĜ�=��#��h����GU|�韺om#�sC���LN�nj�k���,�������=��x��ʏ�~
�^������q�*���e�O���������r�q�*�x�uG��"�q�8$�$�7�1<l�������+������\����	�A�~�����{랇v�����)���吝��}�����7�[����o(����</~�����6U<�4y}^O������߷�37�t�??��sf�߉����ݾX�)�>��S�C��c|��-V~�_�pO��	4r���ŌN��7�~����E����<}�k���E-�
����/�~&�˿%�s��K����V��>(���0vblY>IX}�]��~ȡ�Ρ�o�����'��w��fy&�����W���������@�_�ي��T��U}��Cp}8u��gI��]�������C���!����#|(�c�?�?���<�<��z�~��5��y���x��Y�./^���������o��دA~t�ͱ:.�W���X��w%��T�yq���p����⦻���F�����T~/�:�����.n��8�5͝��3���o�W)�����;��u�\�y]����E�ob�g�JY>$u���Z�V�r��{J��b������/��;S��b���sqz>���}��ϓ�B��B�l,�O��H}��s�_��v����(r>�8\�8����w5/\oh^�����	q�	���:9W>�-~�v�ZGP�ؖ�����s��
������d~�ޤ~���_�ro�ρW~��o���G�~��;�dq�i�O3�_r���Y~w�UM����*��`��b�k���s���y�2�qQ��m͇�]V'�O�o�W{������Ɵk��6��$����g��G���~���������/���D�z~ݹ�L�_��������1��9��zH/]g��x��Uzz�1��%I}��JW�N��!���Z�=��k>F��Ky�c����	V���c{��_����Vy����$�~�֍p~g|^���pV���|�������>�/V��^���[�P�3�3���M��q�K��a�T�]��ً����S~?F�g�խ�i����T����sgU��39�����9;�m=�V��_�.(�������BF���}�^�>�?���}g��������U�<��58>�;zk���R�O�����%�B^��+��s����
�/��st+V�\��U���M^� 6����m	�(�ڍ�>�9J8�q�\e���6��\7�z��^�gc<���O�~z~o��˴SG"��s��s������y��U�Z�qU�h�m�����u��<����T����z���V��Y�o\g�c�W�"�q����}�����������v�����>O�_�?�W:9V������95�|�uq9�3�^/�8t�	߯���v��G����8{/���B��r�������.���׃�=-��:9Q8��1�|�b[-��}V�D�9c]O��޼3�X0���c�Ͼ���!��q�j��?���}X���:eS�����{2�$���<b���"��6��	��}	���������q����6�{��>�����KZ��]��>B����=q'�wb�[xYl��B'����ļ8 ���T���i����������Kc����w;�*.�y�\�-��?��i�|��|a���_n����;B�cԄ#�9��G��9��u�Q������\��<!�!�������UN�?��}6��n�����Mϟ�'R_��W�;���[���F��������*��6\�<���	�Rٯ*>��?��q*��=���W��Q���O��J��9�i�#�~��7�g�]�]��ω�F�v2�GQ��rsq��vw�Wz`���Ɵ�~����ɺ��z~�wٺ�龎�Sl�`��e>jpū�����)Ke���������o�� ��)	=��S�݁�|,���A�ۀ�@|5�����I�����kt}M{�7w
|+v��s�~��/T���2׿���ڟ����%������v��Ιf|>-�����}@���>�E����WP����o�x����o���̙_S���O/�W�-,��H��{r8/N�y����qW?P��;ao�}L�n-����}z^"e!
��ݥ�I?�V��3;v�h����U|�#����ɲ��g�ڊa�@�����޹Q�̡S�g�����3���_u^����y��{��2v��R�_3��ϛT��պ�q'ȳ��N�u>��!^������oj]��!��%��h�Ǐ�#����{�<?B����'��@��b�}ꗇX��:-�_��aN�������߫Ӯ������X}�,��8�}d���c�{@(>���5��U��m��q��u�L��Σ�ϯ��� �sL���gX���'8o����6�y���ϐ�CI�j�5"ߏs}����������ǅ�O�SՓ/�c�e���k��y��L>���W)k���*���)�P��'��8�9e�[f��]�Ǽ��{d�G�p���T��p���s=�slJ�_�_���/�.i���� ���MT��O��8��o��y��W,��{غ�����=/���o<'�}��pgҮ�W��+������sg'	���z��c�s�������N7���<���b*:�4���G\�r�#����O�=g���o����ǐ�@��^_��p���{��������@�����_w�O�~5��x�b���.�u_�Υ~f{D,�*�gĎo�����p���)�r���kU�Q�?�����̔�;�o?m��"Vϛ�oV>s������������ֿГ���]�|QC��⨯/������T~��um�l�M��_���b������:����^���x������b��5ͫ��+�]���<6��"���TyG��p�x�8�s�v��C����' �s8i7��^����������*|�>
���cu�����*�̫�=�A���q�Z���꼨�Ū���ޟac�/p�K!7�����wK�_�D�>&�4����O���9T���"ߗ���?W�ӯ�<�uڃ|������Ǽ��T�b��?����#�����|�R��u^��7X\>�K�saݧ����Es��<�.��	�߯�xg���>8�b'N�~��y��{����=�C��@�/��I��)���N��~^��:���wa�>釼݁/������?�G��S��e�U�6�X�Z��S���T�����������?8���MmH����3#6e\6�����8����Cg�~�x�ʡ��W������|y��ҷ(Y&��E���eq~��x�y��zGҮ�w�����1�C�ݯV9�c�Y\#g�-1����}.«�(�����~_"��,w&x|^�n��kc��>��O5���+��C�]��/F��07/���Y�l���p_��.#F������{�������E������(�IآG	����c��7���O���W��yG��?�C�%��4�p��7vr����6	r�Ƃ����S#�'Ū���ѸҜ��k���v��s����&ϋ�'V���}�p�sF{��E1~/s[#l�?�-����_��x}]��Z���/N�|��a��|��j�ɜx/��m���ށL�ހ_��1ܱ���]�s���?_�y��h���y����{��5���2���8�]�|��Q;���_�'3����Ӊ�����������>g�A��U���{oX�n2����3��������u������H�3���Ξ�g����SX\N�����lߐ�fz#���y��������[��1�K�~%��K�j��������:�Jge7����c�ϯ�����:�W�A�)���\��;���?_�}<*س�|�J�����Y�|�{�k�	�	�9����B�ꡑ��|��� m�|t�,�yX��e�����{J��z<�y,�4<�8j�go��;��n��������7��nZ�(_��<�ۅ��G�@��s�S�g��S����׭kT/��{_�~���>��v�/���WP��E�>_*9$��#�)>����^��;ڛ���9 ���C�\��V��.���~��V�5�r��Pz�(�;�߱X�'A�c�W�߁oG�����/��}i����;�ő��u林��'xܾ��^�a��33׿�|�*N��M�W�W��p;����Z_����],s�$�����ߟ��8�zռ��r^�]C�>+����&>��#�w?`ܟ-p����A��������>��/Ί�%�=����^�׿|���xy{�����1�q=w�	�-K}��k1�[�i��h|�^���?6���U8�@~���^�-Vq���Ϫ�8��Gu�y��/���w�=?svV�GL�i̽g�z�l�?�??(�rżkʘۋ�}��ި�!��|��U��<I�O�}���=����9��S��78a�O�s���^z�II�Xǝ �C���3���Å���*���1�x�|������m+x��q�.�n�u����cv��w9���&t^ix*�W�_r�����Or�:�~o��{����-�F�"������.�T�W���S�yD<�Q�'1��p���x�y�J�t��p�����?COh���������<x�t�������=0����jI?c:Z�>�����G;F���|n��UU�Z����d�9�uz����)���|,�==�ag�؎\(��=W��s\�1O�躏��b��w��/���z���lq�,��=m�[|J����+>���9ķ��4ި|�v����x~�Nߏ#�G^�ע���|����3��ʷ7�C�����������9�C<��������۩<��c8g�zNBg������#���`^d�����x�űj��_�'��q������K
<~^[���}�K�/���^r��A�nI�W|v<�d�twŰ��	��U|8�c8�!?�<^_�S��7Q�����Ɔ���X��O���|>Gx�����ؾT��#N��b�W�bF�s;-3��9�#����wX|��g|�1�O�?�k���k������C?���5�Q}��d6������"��ܯv?s�����_-�s�)���:kG=T��Rn�z@�����3W����.���y�a���֯bGV����X���!�����ʎ+8��ݪ�"�S����\<������~�u��'cO{m7$���zG�����@t�����Wt;9������|��_���O��<+�dJo���~��_�z�&���T%?�˒��n����<~�q<}_a�gǯq{�O��~O�T�����^������Jj�㧝,��\x�?�)��|1�\�S�}��;w�����c�w��ʲN�~K�z�ű:�������g����j+�}���gx澏X��~�ߣ��_�v��c�����}���տ�o�c����m��|�7�#:���~���~#�|Kl�!_d���Wu�����	���O�����R�-Q�@R�`����}�_�i׭�uD��u1>G�І�'���6N|+v�m���<%�R��xчb�����·�_����/�t�U~>��k�#W�:Eq(�C����ˑ^�A������u璌���_��}�Ez���^��U_�����KD�ƣ���<���7���և�:����?�}d�9a\TN�_ ��z�z���ϋ��U���"&�5�Ӌ�j�ڦ�5ΐ�8�(��aY�埥��U��I1�Cu��؉M8�j?��C<ߌ��GS���1}����s��O���۞��y�I����`?���o���x�wŰ��+�*����|�k�����dqC1�7'�Vv�����N����sQ_�q�Z_p�������gȣʏ�39�|i�<p�����	s�+����='��U|;^�w��<�/��y
�	�6g)��E�9�h�3�Ù�'��\-�S����c���u��x,�~���
O���("�sL����;������պ�����U낅�5�'��;��(\��{������*?J������������.�����1~���g��߈�.�x���8�
��u[l@����tX����u��G������n�Ɲ��C�q������?�o?;i�E��gb,o�|n���,U^��)�A7>,��@��M.���yp��G��s��-J?�:�卲1%�|��F�%���O���T�?h_3z*<U E�a�W���Y|���V{,�m~�7bUN��i���1��"����Z�3��O�؞R��}�Ď߶U������L+���1����ڧ9r[����*y�����^f�Ѧ�S�^�����ѽz^�vp�:N�ӏ_Dn7���x�<+�� Y���T�jʏ�/���R7��sy|;[?���ͭ*����{&���O*�P���g�k����O������W���^���[I�������9���s�O`q>@V��e��P������&�$��z�ѱ}���$�]~��gغG�*?�|ܖ���S����?�����:�}�s/z�?W�ie�����T���!�Y���n��/�����|}��?\L�s���~��������m���_�iy���}�a,�	����<e�oqW��0��^�c�י?v ���Z{�M^s�B��]��Vd�p���~7����!w���ٚA?�>-���ޢ>�	ޜ-p�W\��x� ��8)����|]>��I�=�{C��M�>����ks��9����f������*��X�տ�T�%�6�Ž����$x<�e��۳�k�ϣ3�n��<��d}����Y�o���O��_��9��?���������2zN������p��i]����bx�o��_���ю�{�P��1?�W����]�ѡ޶l��}e�!����d&羞%lN�_�OV�"�y�z>������x2�MT��f�+J}^կ�д(?�WT٣��d���;�>�����#�n��cz\�χ�X~�bG��޶f/�9�u%�9l��OM��,������߫�5�����sC����Y��� '����c��ڶ�G�g�ֳ.?�o�����8�?ܟ���iω�w��������u_���m�x?��~K��Ւ���\�<ϡ���%x܎L�����[}�����+�Yܯ�����'�?=wɼLϣ�����������ڻ�?g�X>�(=�>�꽫JO�S�g��Pԟc�����?���L�o�x���,Ζ��2:I�R��s������X]_T�\,�W�=�A�H�W���ท��N�M�#�|�{\����V�A۽=��:j��7��T~)��{z���\�5t�x�{�2y����_�:��	��zF��K�f�s��0מV��08��?���u��O��G�+)�)?�G��u~��y>:���D�\�i�T~�#:쏣��1��s�iVq9�%�o��������<̽�c��<Kv/���Z�:?�z^�W�w1n�1��N���e�އpy����s�x)�q�������sQ�W��T�L:�u�:~f���w�~,�sXW�ا�<;���������U^��qaq�d�O~����7;�t����yrQ�q.�+�]�P�!_�v�Cv��X\��?�?򼬈���d�x>ϔ�^��u��+:Y��<��/������ڊ�=�Z��Ǧ֡�.��&�������c'�Y�T�*���{w?C|�ѹ��ً���A��O�?���oT?�|��Qe_*y��[���x�x}���W�kБ�;�8�W����ņ�����U�-O��W<U��O���ǥ�����}���n��W��}&�w���fx��7��e����]#�D���ߜ�k:נr����_�"��S����j�I/i`��x_R��[F�e�e��j�>��k��
�g���xfE��sN�c~iBOO�փ_�������z4m
��+`{>_*:��+y�ߟ��[�}D>	��8���<�����eݾ��y�����/����'�g�V��1�n�G�}=�9;�(h�</]�3���e��FU�U�0>�A?�9�6�6����s��"�s���&�>D�o��5���Z���ߒ���廊�͍�U���t8t��/���]y�����yL���=�.hޑ�;�
<�?w�X�3��n?����~_����Y�۩�����_Ü�|�s��j�#�_�S,U���'F巰��s^��$Γ��A��y*�u�%��W�0x����,>_��'��I�ϋ����~h��s��w6����$�e�w^A���Ͻݻb����O�u�b<.엟�R:�������8��?CK�!"/d�9��W۟����V��x$�r���B�Y�Y�8�Ic�ȟ����3�0��S�ڭ��3c�R��Y�ll��]`�i^qu���5��w}Ok�ǈ55����+�e���߅1�=|^�>���a����y��ꞓ9�,�Kܟ��G�y��χc�˳�/�+���/�:V�ϾN$��s�s�2�X�q]��/:ڟ_�=���ҟ����+�P�U�Y��0�E~Ύ�f����X6}������S�ݟ�8oS���U>W�)�(���#��w���^`�����b������ӽ>r}����W5yE��m1~�gu��y���h�����K;�1�g�?�����o�ϟkp�����L���.��!7�	��}en��	M�:9�x�L�'ctn�p�k�;z�Z��~�Vy�d��'MS���s�������@�����������ѿ{H�֛n�|��g��7<^���֨���ey���g�}j��V����v�~Q���Gi���Ӧ�3���;�}��������<���9�j�+��~�������V絝�j��=��T�,μ.3��꾅*���K����W�,�_�ײ<�*g>m�\��Q�j�}kk�O�h�$�+�����~M�����ͣ㓌1�>��Ѿ�/��[��j�_e�͙tV�Ό��N�g\�Z����'����]�gb|1ס��^,��;qt�W�υ�1~�(��*�~�2vdvs¾���������;U������L�+�H�ȉ��x�M��E]o��*������r���<�'��\�18O����*�ż7�sH�mM��{��އw�XN�_�S�+m��O��޳�=V(�>��?Y`���mo�~���w�P����Y��)��R��R�α�5�%��U1��S�������WR�9��>˳���s�=�ؕ�u�Q�<������m>�?#��x���@�}���6^�g��,p]wD�g]\=�K�}��_�7��:�P����/�����d=������`_�?����l�{Z���|�9�J����z�c�r� ��p���r���y��W����#d{<�{�9��,믮�?����Sz�����c�<��C"?�{<���>dvj�����J�qQ�O�����8�����|�v_�aۯL�?U��Q<��������T��/�G�3dJ�w���s>㎸3?��M��>��3�o�2��1����O���F\�u�*畟���M�k���_�z<�>�COp��r��[��d�+������_�pw�n�7�W���X}�}�U|�|ĸ<<�?�����i���{�������g2?��[|��hk�y��g�O�d�:��m	�*��گ\�oպ^�gи(�k��������;n<s�?[1���CW�̃�<n���Jk6��޵@8�+�Š�����=��3,��g��Oj�l}[�|cѻ�(���s΂�>���L����?�����m�o��{Y<�M=��N����u���ɛ��KU�������_v�ˡː��=����\����*?����N�<k���+����o��==�;�_Q�������5O)����|[1�'|3�����E�����gq;����-���1ج�v����q�{�����չ?؋߉���Z�Gz]�[����8��D8����G�zY�pv�@�?}�ߟ7c��-U5�\=��������~��F��T��svn��G�3�Z���^��Ok�J'���_����@_��^*�q_�oښi����X��z��]�9ܕ�����C�=�U����w�GT��r���gUx�<T�8�%���K�'��9�u��
��V����!�?���Q����=	�|��_�묘��d��ۦ��x��Ķ��� +�xF����8��T}�'��s/Ѻ��'���v��?�ݗ��~1��~�����"��CĘ|+恿��>h��m��������W�?R�5��-�\�������,ΐ�1�����_+�~Jo4.����/�i��=�ߨ�*;�p�{��i�boQq����ٽ�<8�+?�h��7�G�9`o�A�t?]�K���1�I�g.�>�{u�CR���cD�?��)'�>�O���?��X��-�懟'��&�M~��{�������]�y9h�,��)��r��0��q\S�Q��
���֛>�B��u��+���k�?���'�*��p���`��E}����w>�|��,s���8f�̼�V�.�_���O��Kٝ���1�4��z@�o�?�>�9��,.����>�H��`�0�}�}κ,�v�����V��r��v��A����Gmg+?�}��x�������q��J��R_��4?�˧˹�g��2;5g��'c�unk_���o\�9�����Nߧ	��\�5�<���'b8����Z7x�'/$μ� 7�R���ݹ���w�v��Wx2��څ�C��Wu������9ܟo�|=�qE��)\�M��ap-�|_��p���t���*�D{Q�K��g�'�|Q:��Y(�ֳ���W�nj=��N)\��l�S��D��;�yu���?\?~�կ���(�,���Un�}�?��!�k����qo�����Lȃ�m��]R6�N��2��
��*��ﱜڿ���j�vݾ��������T�m�݌�~�g|]���N�}��{w�>=Z�3�}�Y^��mh|����uI�U|���U��Om��6s�g�{�?z^L��Y���i�8K��+�������Y��6<.�������Lڝ���b[���&�ٷ��R|ܗ���co�����[��~��>�	�Gy����N?�\��w{����������N��Xǹ���zi���;��>�=/��Գ~.���7�lߟ���9h=���k�r�Uz���*^���y@��+�����c�[�/����=�?��������ON�u��=��{dL��=��Wz��ѣ:��#�W��Mk��}��a|��7���s�w�F?i��������L��X�����.�G�����ǋv��|���xg���~�=����c��I�*���Y��k��:�(���>����I+�O����B�s�w:.�Ǣ��#v�{I8bG�`�i�����{�|l��\u������֍�;O��֥&�'}_�g�3�����uj��������M*=�U�E�0>h�|�?�<҇Z}�+_'���c��W~���a>�Y�qOv���֥F��f_��z����F�Gbg_�������Ƈ�uʺ��W�V�\�a<3�a�?�~��+>Ӿ�z#�rf��G����$p�~V�꟩����T���f�g����hܣ���嵱����ޞ����~�\�o<����V���N�e�{O�S�3>��I���&p烖�U����R���\n�	=��,��^����;��{�2��׳�<B^w�U����X�s�e�W��COk�����ߍ�c�mOL�{�Z���pn�%������< ����������Ï��y�r$��rj���	�v]��;��{z��l��t���3����Q��V�+�K
/���uC�o��[ڴ�<�{[�YT�,��E�d����=ⷷ�0&�/M�	�}����<~���\M�/-*oz./�����.��:�I�^��+_]��~C��
�M���=:��[�ƽ���?��}���7�ߙ��/;���.@��n����g�+���<�g�I��P̋�T����	��G�RF��_|r�����9����1�>>l�OOڝ�/��p�K���1�;zo��M��o�y���x��_�c���V�-��;�=9�z���!�����/}����N;���*��9���Nϕ�mm͠�����
P�]ex�� ��������~5�H�o�==o[��X�Nܳ���^�/�!�;��!�կ�?+;��؉Ik^��z�s*��?�ʫ���c,W��%|��g��i[1��x�<��T�k��Oű7��?�~�֯�9U�_���Z?��(�=G��w���c��7�s��h���?2Ə��mr?ָ>�c�)�%��k��yt���.�]k\���(�9ׅ<A�NI�T���58K�Q�)��?W�uDQ�Ͻ�z�=��'p����Z���w�C_��'���q��R�7���7�4�]�w�u
�jv�0q(?���Ӿ��xT�����k��>+��H��9ôSz^�%�u1w?G����U��9�����G��<m|�#��=;����^�u ���ù�����f��5��aΫ�"���u�6���j%�
�93�_=uJR����F���7t�/��x���y�33�Q.K���R��e�Ÿ=/���)�N�Av_��G�s�o4�f�[�5�^��[�U<:s�o�;�c@<�Z�s����|��W��E������*@���mŏ�xqǭ�<���KQ>���N�K�z��1�׎�Z����8!�1������׫�c޹]����d�O�|�u��L�5�]1����a��4���S��{���PTx<O��[(���U�Ū8�&��b�wo����;��_�aX�xKF����O�/1�C:�|��|}w~#���3���??����o׷\�a�.�/���γgq�o�Z����m�g���U9�����Αe�tn�.b�<շ���з���˄?������E_-��~�~������Rű�_�旮��O����G�l�p�g@>�b|/.��9�y�F<�}�Z<�8�]�����h��-�>iw��[��p����o���X�H�g�� /<U�T����*l篵�������}y�~���%���CE3{Dy�\�#i�֏U|�� �*�����w=���Z��!\�پ[e���8��Q��R_��*^G�>����p��C��K껟I��>L�gT�u��������e�k��_�֟���~���e�����H������T�0����������������_�=B���۶�w<>�7ǐ����1��U<�?L=\��H�߯�������y�����,�>��U.�m�S�
4��z/��Y��=��rn��k�����(�cNXfw"�zu*���uzg��c����������E������8.�[zGl�͍�K}��(�M�3��+��!�X����^�'߲�]��&�C6_�u���[}ꟳbw������\���;s �x�׿=�w0`Na�n�_7�N����|9"��c_�<7�����#���W�y*o1��3�[�Y�q
���,�>q���ßh��(�{�C��X�3}��(���������Q��,U���iO��.������A��s;y+Stj[ϓ��"��Mٵ�
8���9y��������U~m�3"__�m���]y^n����Y�}���+�Ӽ��?���7�Ϝ�'���Ľ ̛����[�p�Cv�}�w����՘�9�7�O�5��4���Y���نs�y���s[��}��&��y��w7��J�;����T�U���G�N#����)\�P��5|�{=��_ʃ�WV���w��|�(�qN��,n���n� S[���c��>�1���A�q�_ᬧ�3�q~�wE����>��o����/��]cy{P�����P�>;r{zV���Syn��=��|tyS�hN�j�W+<ӫ��cu^�ZG����q�����������s��L��{���dB�����w;gJ�8�jN�����D��O�ֿn/����u��g�Q��@����������yN���˕�P�;�y�q�zB����A���b��{����F��x�n�9'n�e��U���#V�yi�6�H��=)r?��'���Kz�꫿��S�y�7�;y=nG�?#�q��X�����H� G���w]|u�|Q���S���g�9�L��~~W�G��OW��p��*�i����_�����N󈖽����2'.D����,����x��=�?=�<5��ߖ�w�*����oB}]/뾒���<X��)��R�m��X�o�~>֛��?Y������p�ٷ���x�������v?�>E�:��O�m���Vr�y��X=W[�OT�͙�z�a���L���ӌ�������S�g]GT��U��|{v�ó��[
\��S<�ü����\��������v���c	��řQ��7�9�Sߓ���4�	<���ʛ�뒝���U��zI��f�Z��L����a��}����kFO%�>O���Ѹw�7�[�3��x�#�_�a.���U�C�/Ƨ�G���OX4��~}C��N�sF���y~����I�?n$b��b��'%���̯�/�gt�f��;�W�	.'޶�;�H'>��3�_���b}�ϝ�L��y۰�N�=�G"�'�s�������=�#>.�Q��u����]�f�ۺ�n�����m�\A^����+�#�@��?~O�[�fx��u��aq�5�k�=����J��*�1���aݏ8�s}���q�\O�?��2���aM�����[�T�Ff~�"V׳�M��|W��9�s���K�����w�p���s���b���>�������Q��,��ί���D���Jϔ���y�ؑ�'$�}~���fv��s��=���B���c��Q�_�G�w�.�c����}k���q�����Ƿ&x\���1���S�q==����(��1o}J��ݞ��k��K5�s㽕?\�yx�R�W��{����w(<��y�=9��9��\��9 �ez��L�Y�V�e�T���z�����oGc�#a�4��`.f�*>|���}���<C��b�W�e�8�Ңp���D���_N�`������]�[�����a��D����?ۘ��4���U�B�?{�>�ac9<G�Z��^|u�X> �_�k�y �W�1kw��2��������c�}���w$�����3�'�>r��}4�_���^W������7�X�u]��ό�2'�G9��r:�#��v�/��:ytG��.�8��ݱ�Z<.��C_#;��.�����~����ۘ����g��e��ʾ/~cq�G����v���~��;�c��ՙ�����x��)}X�3�����*�EY
��D�șI�u~ԙ	|O�q�#��a�������ej~M���1C�܎G�$����V��{���5��m"F���Գ7F��?��[��\�x�SK���g��eSv�:$��*?<�����&�k���w�'��Z2����q9h�9Y���x�N�����T��Z�]E���H������ZM���zs��\��پo��eY��;^�~��������v��z��m���I���8)n����������R��X���|�J/�m�;b����y����O�[1g������<��xZ�{PR�������s��vf���-��k"?���I����[�/}bo��~,|=�5���ȼ�������m,}WR�駝����9~��\<��T�0.w����s�4.wiR�۝��e��Yy��Sqi�㐍������~;���b���u~o�}����8�FQ4_��?����7��y��<�*>��	�Qܯ�y�{�x�w���?�]�}������;�X�U��*�2I8�H�~�VC�ؼ�_/~���i�ھo��w����=���{�z������F�'h}�;�d���<�[�}\�?�=s�^0�;ľ�	�3������)�zrƠ_��̽�s�#���.X,����o�\@���j���/��V鍭�L�:��V��U��΍_��6������u��9y���/�z?T�������ݟ��{�{��P�,���i����'�4��������	膓b��X�/�U�8.w���\��q��K�WT��F��x����IO[L������Ƚ�?
F�S,���������?4r���wcL2}B^drX����R����d~��S��Sz�w�؟��ap-_��~6���ϗ��y�u�A�x�����/���ʯ֢���^������⹺�7c,W������X>��e��c��^�~�����s�-�_�tW��9=,�_i���{��Ԏ��_�~?�׃�~�iJN�/��zoRu�����o���͗ϕ�M٩*>�`J�O��㐧p�_���+?��_���	��qu�c3ry�W���7���ֿK�C��X��V�����I�N�b^k��:��0�sj���}X���_�����w��1�ϼ0���u�^I�j�E������ٟ�}�ώ��xV_�З�����uМ{bU�x~f���o
����!��Īߢej�P�g��ex*��ϫ�O�Y1����;�0V���^�M8�ӷb<�{�?5�T8��}��'�>��~�}n�Ͳ�>�b��2�����,.�gu��"O�X姯˪x/�:}>GON�g���㹫��|��}�A��-�U�^���1����M�gh'~��3�1.�~P�>B�x�v�w_����A����^#�+ڔL>����-ď�U�M��7�R���#��[%'U|���܃�#��;T�����g��]g]�a��x���8+����\6��"�/�� =������}Z*}�v�v����s��k�o���9k�!�O���S��~#�S�q��x�S9�;��.�sZ���;k��o�y�u�eQǣ�q��o>�7�g؝,���(�a}>�&����5��T�������?������g�X?T�j�B6_�~�_�%V�j?���*�������O���6����Y*z��������\���*�S9���a���g+�_����WoO�c�k����;����C;��g�?�����ę��u�8-������:�o�g29!Ms��S������Z��f�%7���o��T����C����vo�p�e����}
���[���z��������[�;��ל����9*�3�o��oq���x~�Ƶ��ս��
��6�>5���X������'��6��Hϲ|N��|[?T�z�R����r�tg��G�������׃�*�;��u	�u��]��8n�yvy���𣨟�V1�/j������9�����Ww�)ϕ=u��M����Ф�~�֧?��D<
{����{�1_0�q��S�yns�������ג����?��]��;��Lï�!+~�K[Ì�#vK���2}�zX��ĵO�/��$_�����W�L�e�β��o
=
�����W�'��� ��qw=3�o]��{�+����8ό\?��s�W��V������h�ޖ�ohS��A�4�������X��Ū���,����X�{�g�x���	=n�G>W�~���2����{f����s|վ'�p��1^����_����u烲~�~��;^�%�P&�Σ�������{�Q�����P��h��H��޷c?|��
<Y>����B��q������g���s�v�<�T��B��N�Z��\�+;�S�C��jq�����@�>���=Y�s�,����4OF���?�Q3蜊��7S�T��n�{Ň��i���ϓ��q;����^��ד����g\?W�
�[}��~��̞�?C�@�u^������ߘ���w��p=���K��>�y;f�3w�}�u#b����z�+���9�vNzվ7��'��ߑ��/��������u?����Q�|�d��|w9�>��U1ܯ��tV�?��ݞ����c��������]�j���3�a���Й��}?�t.�v��gĪ�1~�Q��|X�w^��q`�2�|a��bm���>���C�O]�u*o�t\^�w9�z��w:���^L�G�z��w��Y����w�ԯ�c������h�/O��\O-���|��ڄ�s�ꍽ����w,�ޞc�~�0�m�~��E�*��6��>/�6��~^�~���������a/�:�Ki�p�Ӡ�4���+�iaoo�K�S�)��� �~���ߨ|�;h|`�g�j<���l�zt�8�Ο���<8�@ۉ�_�o�R_�����	��$.���/�{
��X�L��k��*'�q��������q�7�l����ޫ<�O�!�!����j��N��:����x|�e�{�2<��T��K�e4���q��oN<��J��s7��^�o�A_����X�)�:O�� ��A��5����a�o8��ھ+������>Ke/8w2�e����;��u�����%ş�������>V�IC�����y�c�����Z�o5���U��/G��:�H�;�Z�����e��o��*��eo��x��9��Y��4�]f��7�O�ɴ�����!�eʏҒͯ�Ƌ?��9�7�O��ϩ{f"�<O���%�����5�C�'ߩ}D�9��b���q����W��{=�2�߽l`��7E}�˜����CGu�?���u��gE�A���O�����?�U���ǟY/<���2=��/��Z����I�y�h�o|�����m���Yuݼ���,}j��{�7��ٿI�����J�C:�rkϘ[1������ƅ�]��w�x��:�߫����<5��<�y�08����v~�(����_�sU�xxy����X�[ş]��ˀ�,�$p��Ü��v9a�2i�j�u���,.�X�ι�ʓ��c�ϳ<.��j���u��T���n5_�T~��N~�9�}���~m�����RO�s�";H�[���1�_�������2��]���v����\�\T���U����?����g6�������/��!�gV/�A�ҟ�Y��#�y3��E�ű;�03~[�����3΂|c��C5.��$J?����ɓ��C������L��ܟ] o�bȳ�@��9y2�ſ�9���>Y�`��Ƶ��ˈ'�OD�g�gu����g~���~�g
����xTz����W���x9��׌����N���z�������~����Nٝ���Ƀ%�s�i�����{�Ӈ�b�w<����]�{��<��A;��[�S��>�&�}��a_Q��=�+c�|�o���c����Ư�o(����������|�O�'��yt�?%��U���p�Q2>xܒ������#_�/���[���3��+����p%���۬�؈;�f��u7>.0V�}#�,V�+^��c-�;��%p�������S��G����sQ�gG=I[5WoW����|~��U|{#����ɭ�?���|��������W���f��g��|Y<b�o����:=����_g�U/-��*����$����&��k��w���s'�,�Q��j]��c�z�����ޤ���v)�d��Ω��uvA�-�x��x��ÑK�qB��`����G�����+0���c�zp�߫��$J��yk��������E>n�r 9:��q�3�o��k��}s<U�%�[;eg�\�������w��R?���O8'��gy^"��y��z�����qip��"��x��M��� .ǃ���w���n���N�[G6��/=ߺ�}:�֢݊�r>���~�~�����S �}D���&V�6��_�m�^g����s��z�%�v{;�_=_�|�gT�̑�l������5������;7^T鷊�o7��}��/�d|��	�����U>�'�Y�������G�����&��_�X�;z��U��3�|g�8��~�
���g�#~"u�����r�u����zzߕ��9�Q�E����n�F��
�:��w�nF�����T�$�q���_Q�OF���Cb'����R�hB���V���v�g�_��?��T�(����w�]�s��E�5�{�x��ע�H:��G����P�<�;��U��nG*�A9?v|e���<�������k��T�D����5�ex?���@�ev�ϡf�R�����������t��[N�U|�� �aN|T�[����ݗ��|r�s���������\Of��;������wK�?���>������8�����S������2�n�|���7�X�k#�7���cF���g�a�oU����ӫ�Q�U�H�WvAK�WT���c�����/��I�@~��/�pإK~��P�K�����Yܲ��@>��<��U|��<dqK߇��z��tcR��_����>��댘g��>	Ʋ	������m����������S��y��ǀΆ�%V�m#�s�/�G_w���h>h{Q�;�|�Guo��a���[���C5��}����x��7���N�I�:�>8=,�<��� ����O�W�=�pS��^��1m����[[�M��\���.@����Wƪ]^Ī?��u��ٔg�ϫ:�K�/�������~�I1��j|I۝�S��B�n�y�zO��;{h�'��[}�2����i�m<�u]�y�����uDE��9/�y���0���?�Ϻ-���5mw��3,����w�M߯�p���1��c׼=��*�S�W8�T�;���ڼ)=��;'%�t������<����־0�{p{��n����̱�,>���o��n�A� �'��N#�u5L������@�����~�}w��}U��W�7��(��V�Z{|@�����dY���p�#�Oz}�j|���F�K*��\���y]���w��#��k[���U�d�_�~N���<�����>N%�����$?1�)�����;7^4��x}�Y�`?<�_�G��v�=�.�C�\¡3`��}����cOu�Vv��z������t�7�/��۹¿����TrH:�W�wt�~:aټp;�Fy�<�H�,�/�+���*��p���'��ۓb�`]���HG:�q������X*=�6�vU?/;�躛�riB'�@�s����X��3���tp_f�cgfvS����þ,�3`��uy���=�����	�g���!�;>^[��C�zfi�!�+b�)�S}X��7��bY�s�d���嵮ҩ�er��7;��G����˳��Ù?vo���'�l趫w�������0�/�5���X������O�������j���c���܏����Yu6��G�~²q������G\(�����J�2�����}1}������{�kixN��X��kTţ*;���y{��U/	���q�;�X��x{�j�k��+���s��5����qe�wU�T��ݞ2�
��
�߻׵�����st�_����{pGj��_T����B�s/�0��_`��{�}����E�@�����[��N}����S��G.?���],��+X$��'��,Urş9���j|���/8�{P!���V��ŭ��y�}�;�+��#���|B�[�G��X�'��oEu_���q���7�g�ߥ��u�{J��/����~������~9�/��w�}��[�7��Xoݹ�j3x6.�v��/��j=��3�|�9b�_������5�?w��z~W��y�������pl��;�w
�s:.���U�(/�x�)	��dO������3�O�X|�5��t���9q��1�o|��������y�ur>G���E��������X��h������?Y�E5���y r{�x΍���G	q���A/�U�{�����l��������j^�f��'�<%_W~8�s����עx��K�Γt>s�r,V�<�ܥQ�/�_�K���c�?�;�r��O￁ϛ�;�?ְ��3��co}��o��}V��g��ܧ>l����&���~(b�y��1������]r;W�
�_}sQ�m����-��}����C.p�*r�t�����*������$��Z���,>�Sy�Y��w���k���N���d]�z��e1������EQǩT��B1^G����)�����LO��w~�T8�)�2���c����U�Ǘ�s�J��z��q.����K]?޻ӎ\��w��}���O�_����{�}��~M�#||��.-�����t:ٞ��ur�n�������E�yd�����o����Y�R=�31ĵ�Ͽ���::�kb������o�+9�|���m��5�<�`��s����|���ύ��IV�%���������W�ߑ����F�����x�~n�7�����g�K)�����o���/�!�N���b>r���������d������K��/���w�،al?����[��j4oj�z�q/�S�����ޯ�v�cA8��K{��.`?�ޫ����܉,>�c;��ҧ��Y�:��񫞡^zDQ���w����)�����s�`���38|��q���u��l}T��Jߺ��;��~K��D=��ou8�֝�����D��8���������]X�X�����W��3��������u_���s�`�,���_]�W�<�Î�p7����ن�'���|�cU��^��+���ʟ�{��~f��o���U�F����۸A5/6�~/��x76��s��E��k������@~��g�p����<�~��xiQ>�C�/�o�������M�W�ui�q��~���=�;�������>a֯9��X�_�����XkJ�ǡ��ǐ��3c�P���U���V��qW�6w�Q���������+z|��}r���ގ�瘪{c�ݩs���?c�YߣD�Ī?�3�E~=���&�����z�&tV���~���U>?����X=�}ME�h3�����ֿ���?��b��g��n�4oG�z?Xv.`_���������������ɷ����^�������US�T��z/�n��*ߌ���'�/�������㮝_�T�e���:?P�6R���*��hp������7��T�q�.��6ن����m�Ϛ��M��l{���9�3�?�g��=�q�����k\�`��d\��˜8���fݎ�^�ԯ��<=�����u�]�߻�躣��8G���Q��0V��_���m¾��,~ޓ�X�g��7�_�ω!'���v]��qݏ�u�>���y���߫y�[���V���������c�"=��_ů��^�zi_���������s�^W}���,�D���{����.�����*���xS���cY�*>�}$=��l����2������0�f}a��&�QT�1���|�9�����fX;S~�u�q<'bC�皤��y�U����6�3^������ء�9�׫�	�.8'�Y����Y����9�g��`j���P��:/�;{&�L�x�����;�{:���'V�k�������TI���|�l�*���[ݓ�?�������N{�������C`���w��ע���2w�P�?
��\���W�.�/*'|ʞ��ѯ򌽸�C,�c�*��{�g���g��8�|��{v��>m�u*��O�U����ڵe��|��Tq���a�q�:T�sꓞ�Θ\ծ����;�����v�~��EBϱ�];)��q�?��j��������f
���v��:��v��?Ҩx�u�cc,��K��3��}7�7�������&^T���3����#`�U��)���׉s�����x�w���E������/=�Q�j�7��^���y�'�t8�(\�+���!�֭	����{/������yq��OY���xq�>A�kx��=�qC��~���?�هڈܟ$�>�G�L�o�y�,�NQ~*r�w�����(�3Y�k�r�{~n�!��_��s�����E���#�l�}�>�AO��߲�h%��+�k�k_��'�S����Y�Ε�[��6U�_�:�kU�"����#�R��+��������������� ���];�S�l��g�5�]ڗG~�Z{m��`L�Dxha���-�x��xl�4���W�,X\~�'_�����\��O!p������뙪_<�����������92�K껞��s�x�\T�e9ԯ�}�czr�rB�z�ly�;��̯��G����p�����<��Y�Zu���9�����nx��S���1�C��Y�*n��r�W�_��Y\���Y��~0ƅ�f+�Y��}fz��F:����mЅ�����X�g�W���[�;���O&�}�Ҟ4<����o����u{�{J��ana���}���=�����Wz29���~]wg�Ud����2�w����p�u?N�@���1��E�eZ�_�s�Uy����{�*?Y���X�~�,.��5.�����7n������ս>�*�|���oռY]���.��9Ƈ��y��a����V�wL��/oE-�j�pw�w���z��������|s��c�G�v��sR��b��W�8O�w1�^�U��7ǠT�k<ξj�Gi|���?�Qا;�x;r0����g�z�<?���9��Sz������5P[�/�*��>�?Z=��6���o�!ր8�o�x\"vκOѯ�'DR��y��_���8����칶���o��؉��\Uz[��Tv��Tt���ýN�}�����1�ۚ�Y�߅��X�'��g�!��A=g�y��^'��s��t>j���3:�K���1�Ǜ?_���4��{��=��i��~m��b����Xw��2vx�x���|��08�����\��=�_�y�K�I���j�I��[�|V�պC�e:8�����{ܯ£��ٺ�h�ǅ�(3%��,��p�����sU\��	���������;]/8�+�b���v�_/�<#��U������ތ�� |>`����ϋ||O�y��S:n����������>U�ޓ��+|�ۺw�zm�����u���8c>���}��Oλ�b<����>zE��o�q�ѩ��eѮ�Ѣ����#��Τ��_�~ێs5�q��c��z��{{*>P�;*zt�d�۸�g�
���X��g�g��;����sO3zx/���8���ؓ�?�f��9h����)}H��']��of�v���.^������Ww����7��-+�����^ϯ��׷'�׼���h���>��4��$��2C3*ͬ��2(�
Fp�q�&q�@�C��F���cb���Wݳ�﷿�:{�����߹��:�ƪU�ַj�<�����#mH�z��W_W����ܽ8ࣺ8:w�~�SV���/8++�Cח�5�����&K���oZ_�Ͼ��U>'�X��έ�z����\��n >���نƋ��A}��{A>������n����\��5�������ieG�0��g�l�����Ͽ��\gra���w]����u2�[��1|�όO�H����E�tM<�ا���p}�W6ŧ5?&^�5�����Nt���/z�ރ�8U>�^�0�%��kv�:��O,$�C�-���3��[��q�,���t�T��7���&c{�ΡNJ��r�S��G��Z>�w�U�~���@�./����;�[�p�˂�Y\#�ۺ�+����:f�����o�����?Y�)���G�OwN���*v�+��z}䟕��9?W��I�l�+���z����o�����V�H�^��up=5ޯ�P�X��٤�.����Z=�a�S�2ӟ�u�	}����~�+Ϳ�x�!<@��e��ϳ�Жyh����~��E���[D?LtԟzrC׬��s�������|e�K�}.k�߷qg�=�r��[pz���{/���F�����[�4������Wo����Y���?3�wD���9����CfO�}�Q����&�����v���*zN���Y���\^�~���q���S�g3��})��8�c���7tG�Z_�`q�vi�y8��-�m_v�����c���9�G}��q�kݴ/���$?���SF}����$)��bY����� ?�����2>oEx��ڠ�ں�<�������+�3}�}�����ʳ����q��~�������纚�c�rU.��^qyo����p�����J�έZ�Y������ �Ϸ��?������d�9�}����e�ߊ�2�%���N����^����^Sۍ��g�ry�5���)���L��Ş����{���śa�s�>�g]� ~C�b�ԧsj�>S��;��C��2��v����Y�տ�����~�Hz�N�����d/���iA~ƣfv�]x�:��Vz/~�u��������;�D�xzV�V����A|���\�)�!����?��}=j��z����G�Ոϭ���ȧ|�n��:����� ���Z�O����Cj>]�";�p�ה�n�������B~�{�7�I������:p�nq?���C��������������ƧT>�*+�ׇ����t�g�O��v�D�������0Dg�g�'G�������#�O����c��=��2�_V���Ԡ]'$��Bt��Fߪ4���ϱ�x�/�ϗ��#�ОD�-z��|�>g�ә���\��0:�p��Y������c�V�;A�V�G�?Qݠ��;e�'D�j�c�y�󲲵��~�� �|�y��h�Y���)�Y��f����u���w�XV�~CЮ����������j�z���t�"|�X���l}ޕ���~\��?�~��8-��L�3����:^8�8O��XD岼��`��6��\_�#�\�I�{�K���A�_������d��L�"��VF��g��S{�@׹�qEt����i�g�"�=ûȞW�Du���nP������K�N��~*ã~A����ϖ�0N8�����,nS4�u3����1��A�gt�t���o*][p�L��F���r���Q��JTO:�xym�b�ў��cj��/Ex!�Kd���➔_����t���2��|�B�{��~'��l�*NR���ٻ����A�TN��\���8϶q?[�[�������g��5y<7��(?�ҵ�'d�,繝���?�jOXl������~cy��`��%֓]�N�����ɻ�ԟj�G����̯��l�h������@��68"�j��Zwב��j��?�|�"�p5�&�?��2}����/�j���$�A��H� h(��^����Y�x���L����{�:��ʍ��'6�k|�"�ݗ?_��l]���o�օ�<����ַ��A��g��7 ]u��k��蟱���G�8˿)���x_�y��Տ�x�?���������v7��j�=���*��>W�;�'Y\bKl����韖sm���T�-��,�zZZ������)l���8b�������.2�=W���B�`ߓ�3�K{3��Uu^�%{wE'��֧��'��r}u-�tP�Ô���N�ya^�J�f�=��V�orzF����c�����
��z2��~�����G����g|2�1�����O�k��٧6����6O�߲xA�X#��O�)�1������*MuIt_����{��~�!�>^[i����{^XO�3�t�w)@�r�>X�wg]}�_�z�/Ͼ��}���iy���󈃊��l>�<Խ���������W˳���F��/�N&��^|(Ց�+M���y��\�����'e��(�i�Z�o����"�gΟ�+2���c;��`���q��d:��h�3�p��{{5/���>�S%��������S���⼵��UNԇ�2��4��(�'�k3�oe]��"+?��X���[?��2�|�pM�ͧ-���U�t}G;-åd�-[w�*����_�
�emA��7�v����+�K�i�o�v��t=�q�G�&���_�g�O��\b�j���2��y0a�׺�>�~Wͫ������9��v�ߒϳl݂�5>�.dw�N�_`zvnk����5�9	�|n>�O�;�~�=e��~]}6�<�Net�{s�E���<�L��~�T]㚽�|���U�de[Fz�"��Y�ĬPN[���^e�e�N�(���<���şX[!�ޑ9�m�[�x����юm9�t,��'��v_�%��$����2�Kj>�����~;�D�M~a���	�x&/ZO�cc�:�oe\K�U��U�?q�̮�I�~k����wLW�Ey4;C�qxܒ�����R�ז�/+�E���:�)?&l��V���vrƧU��~�c�7��'A?�FtMO">��OQ�&�9(.����i��#���������>G��`�{�����3��k��-V�o�_���MY\e���O�W(/(w_[�Lczb|6nÔ6���G�G^G�qzV�U�?��4�6����ݔ~�x�_�xί��|r�n���~B������@���z�7�����?տj��~��پF}���k�F�YVw�4&���b�1����F���̿Gx���+����"['"���v齕����癄��H�?�8E�#:��>��~{gV�C1����T�7,w�|.�{z�6�j��x|����>K�<f���+	�t�џY��%��+]��]x���+q~�t��`��czCe��_��ex?ӷ�8�������e�Am_�a>��Ω�v�u�����s��?���0���������?P� 1����<��Gи�/�q�LL<o��?�V�o�g�PVO�=�g���lG�M+c�B&���fm����7�/�s���؃�{���Mz�ϵy��L��~���v�i�+�}�ghס�i������sx�0?��g���n��яmx�/�6��/�*~�����/ٺ�~�s���LYŵV�����(G�t���Ϸzd��a=sK��6�{(���ڄ�Z\�Mi��?|_U������C��x�l�;��oݟ�݋�k��W#DǄ|.��'������!����յ�J�\2�����2�g�_�7z��H~�����<���L���E�3�a�c����OT�qM��=�����/��G%��q����Иv��O��d���������Q2֫�]��	_^��?���L.��Y�oy/!ұ�<G[��7�y>��ϯ�r�/�3�{�=z�g��-�G\4��J�5����[�o����u�~���{���~E\����_FW}�/d��D����iD��9�Ϧ'��uI�p=���V����Y�락(^
�O�ϊu<����o���%NE�G���{U�s%޷r�r���̏���!�߰��|�}1��PO����7M|Nj�����Ʉ�{��y3�m�f<O�y"��~)�_�����>�3<?���1�At/&���ԮxP�u��y���3e<����G�~'��F�
�ߚ~�����~P��%�O;_��p�]]��8�L�G�k���/+Y����;�z��z��ҭ?��la�sQ�mw�/+������#I~����g�+$?��q�콩� 2^wL~�?���<2rTO���JS_X>����d�Bv�>�g)V�*���c?�9�e��D?g�G�o��q�foe|�?�>��L�m�L�\��{��[=?L�po�J��{�����hW����D��*~����۬>�����@��_:��VMh�ϓ�g|�yݾ�E^��G$�GlS~�9�m]�v��g���r�o�V��r�����[�S��g?�ѵ�N�3��?��9+��q����'�1;��iz�!D?�~�~{ ���5�ۚ�����q�zΖ��UV{�O/?������!��-2�������%g��iY�n�h���X�WVcR�f��ciC�z@���)3?|�O�zN����(G�*�Kl�X���|��/��H��B���(GH��.KY�g�k=/�ݳʯ���e����<^��}����A�5��5�����������N��X���1�>F��w�������l]��SzI�����l�h~��d<ou�8����cvZ�~����Z��!�_�硎�a��'־+:`�q>U�gV����>u�����g{�X�#��pM�q��r6�����xe�,�s�^�T���)��!��Dz�l���}�LG��uz#�;毲�Y�]O�g�y�{�}�H�[�y�<�@���O�OK<v�j��x�	�_A���1ٟ���Ԥq�P.�N�?�Ӟ'�u�Õ��q��?�8���aH��F<���
�ׇ!d�Xj���#�'�v��'y^5�ڇoL��f�n���QB��ߘO_~�v�Ͳ������'���WT^�?��,�m=��/��`^���b�n~w1���g�U빭�wSt�ˌ�}�~�yA},��mޗY�����������7gx?�֛M��>����q}H羛�3{q!}����f|�"j�%�Ӭ������A�=�ٱ�Χ����I��O�������J�ve��Ō���>�ϣ�����#;�w����3ǹ���_�޸K������3;w����������-{��۳�B��sL��T�������L�@��Ml�v��w<�#��R�)�g��s�L_!��i�ޯaj��sB�} -���e�}{P�����oS�!��́��֩��c|��7/�v�}�d���WR_��^�l?k��?���y�N�^��rh��|�X��#�������Y~K<�ٸ�p}����`���L��{�@�\dt�?Dx���W�-~>�:��k�c��(y�"�7���$>/��"�<���\��Z'�g�{����������;L�̯h�@���#����8{sͷ��f��;A���C���.��&��^+��2�����F���^��!Zw��K#>:>ѽu�<#n�g�/-���?�;po�W���u��Zw<��CV��Un��f�D�������6�}�u�k,J{(�/��3���������n���'�g��=c�r���e~@���(��K��H�u(³��"=�/ۧ�\������ͼ�� ��~�nY�������U^OM~�L�d��ؿ�����Y��ra�g�����O׍K4����h?�MVghO�I~l����pm��:�xl<_��Y����q|��K��O�G���V�)�Ǘ�!Y}6+}���k�·}�>�>����-����/3��_����7���>V����y��z���!�3�=k/��/.�w�ʮ�8�6�u�[�/�������~h�ϩJ;!���2�n]}0?��1��~��sXr=��p �?+��]H�±g��9����l�(�����㸞��R�� ?�|or����[���8���ս��
��z^�z���3��Zj���0����Gj=L�q�#�ׇ��q��X�qQyJ��%��A�ܖ{(f's����f���~0;���_�B��q�7,3j���zX��:e����x\�o���ͱ>H������KqZ�AV�Z���8�zY͝�!��y��例�m��k�e�2��������o�t�c��+��ߩUOfvƵ�u���T�y�A��7���?��"��X?h{q�`�O�����d���\�?����|_�kk�t/���]�6�����+�n���Y�ծ��E�g��;W���h�j,��e|�g�>c&G��_�����R����ϭ�LQ�~y�|S�q}�>T ��<Ň�A�M�uV��?�������{GR.���eeK�ɽ@B��ql=�g���nd��%^_l���
��������(��a2?|4�/���e�g�M�ۉ��B�-���y�x��܌~�>�_��v����|�����ڥ��K1��P��7�7�o[�m�oh�����?�E�y�%��`����\w�
���Xև��q������O����g�yv�ae�ι���cQ=��h\2;�(����E��D~�c\O.���s�Ob����t��������q�5�~��K��X}���7�u����m�O},�c��	��6��OL}�'e�����Jc;��5�?$󇳼ܸ�?;!�|��RL8��4������A��,e��݃�q���f�?�!�G���lߡsI�R����g�ov�T{OA}�9S�E�����@��C��&�.��L���}g�e�7U������r�͓l�e��������7��,G�g��Yw���,�ﴜ˃������h8^<6���t���X.��LV:�֠��?��L�8�%�g��y���:bi�y:�3�Ή����S�َ:Q��w�m6�i��=���m���$�}�O�.nI�W���@t][ʞ`�2�	��j3�9��g�W�$ҮY��Le�{��o�{�Y��w|�)�O嫶��J����q�FM�~3���z�C��y��dv���W�U��i�t����Y��N�˵g[�>�)��k��aJ?��G~0ίq�SV8��|�8���k��]��v�Z1��ߴ���D|�"�7qR�������a��uY����e���׵+d��n���k���>��c��y%��r��2�K]ge^̾5�Ӻ�f�ٓ*G'>�]4ϣyh85�{��_���ɿ+~>�����z¾o�ǲZ��d�~��0�����mz�u�O�2�����[��,ezU����*�_�x��{j5f6ƃ2{�B��*�W�묽���wm��H@:⋰\-��+�B�^S��7����o��<�el/ރ�%��g��z����� ���?.��ri��b%�]4���n�o�?�7�d��Q?���� �_�8��{
Y�H��<Ӌ��P��I�}���P�Eץ�����c���sC�_(�ʑ�Y��%�뀮�I=w?#�8W��u�u㇂rE��l�����D:���ԗ��qI���Y�'���GX�s���OV�,�w�c�S���Z��?�~	�/��ܛzN��rA`���ŗ����]w����g�G2��i4.��_�k)���b�D�[�?*�>�ّ�ъ���ߗ��}�]������������Z~���N���J���FY{1![�7��V����7�y��I�?�s�#���q<�G�Ή��[�}���/���{d�����!���kX.���"����?�w2>��]��5i�]�����w,1.S���u����ܝ�A�#U���2X��w'��~�΃P��=Z��y��$�s?��x=�M���� ���>�%�k-�&wY=����n�o}�: �7���s��ܙ��Yyٸ0ę|�͞��x�zI�T�����ʵ���x�~�~��3���)���b�	�O��d劌�yɷ�w5N��<�K�_���ʞD{>�������7���6Sz＄n��p켞>�|5��.�w��q��?���9S�[�T ������d�������C��'pCm��%�����������xn��Y&�O�;j�?5�)��iџS�*���g��d<�,.����1?!�y�nY��ď;����c�8+����[��y]����_2c���a�_�"����8o����w��i�}y\��ٳsFk[����G{R1Ϭuy�8��lR��w�������<���rw��lύ����j�պ`\k?������2�Բ��g��'�������O���>W��>"~��Y��b귃��f�kߜߟw��ﯟ�ODܔ�ͬߟ��]V.���>Nd,/������O�{�������h�3.1+7�g���=�r��z.�s��>���������d߮�r���~��K�{͸>7 ��!?�FF?S�O�~�P���<�D��u�א�{�";��gv�Z1����8�}��q��Q������<d|�%�kK��bo��U�lq�����Bt�OD��]�{�2���7����*~�=�Z�������@��|����9�g����;e�e�Q}���du~�Q��T���5��@�86���9���Y�g�f���������}"��\�?!��[��g�����������>O�����?�ϛ2�[>Vy��zfz��]��2�Q����t&�ٺ��s^��&��|Db��j�}��ZYٽ�'h�u	����v�8�V�9����m�K|�IVsQ��mI�Q=? c{R��q���k�ii��f�����i���3��������0�'��+��7Q{-��;������w{y�m��H�Ǹ>*������2�C^�����g|���#��n]���X�1���?�op?�=�^��b�Ύ�D�=�;X���K���v��Q��ee[��pm�.�_���ݬϛI=���r-�������c�������Q�
������u�v��s7l/��|�w= �V=f)�+2��~ӊ�����h?D��ϹN���7��$�{�k�eqn�Ս�.,1�,���8�s�r�yU�2<yv�r�s"�sx���'$��~?����c]B�� �#������Q>�.+�ڔ���'�n�����xߧ����#���g򥶽�u���~��U��#2��`|c|���UG��i��#����z)[-'������W�~=���Yt^���L�q�����j~���m{��� ������F7���N�/�s����V��q�xD����lY��yn�p@o�o�d}V[lt�����{�"�8?���Eq�j?<=�'���Y��q��>iio�{G�C:��k'���Wߦ��U�G�����zN�� f�d�(����#��}�b��V�1ZO���x=b�V����ڳB\�ٝ�ړ�NVwx��������?�5��h��~��Uu^�'g�@\"���ql^����p+��繎ￔU��@|��exT{�y�C��6����2<m&��OL���������7�81�q��G��IV�콱\���1�{F֮����qD�a~5��7�2���-ٺ�՟�<����t��뎽o�߇b�v�x;�R�~׬�VW��eo�2����̠�"��X�������;�Y׽3�������HG&���'�[;[�%\�#>��[����8�cn��z���{Qym0��cG��%�>"q��>�:�����C�[l>�:�����Ŀ����T�F�~ےU�+]�v>]Or���������bv�~8)+l���������~�l��u��~"���z#�?���r�_��f{�#\ǣ���1���*;��g�E<�1.�D7�
���������n[_�x���&�%b?d��p��8֫���9⾐n���6-���5���o�eM�C��9���q|>��K�k�����9�o�|��c�жȞ��=�'���S�nW�ވnߝ���V�e�?A|�y��������kK��X3\����d�K��	ճe~��+������}���j,Wyߘ�9J�l��G����H��w��x^��K���^�)�g�ǲu�D}���|A뭲�s���X]�/�v����n��U_�@����I�OV��vK�gl�ُ�����n�%q�����[Z��Gz��v!����'��Gf���7�'�U�U߾�n���b��wK�=���E@G�7�t�>:'�2���3�\�;	}P.��'���3����Zb}e�f����#|��:o����9g8��W9W��������7�%~w��e�,����>:�G�d�qe�?�}��^-��s�Ȟפ���X�����+�>���[/"<�&]۾�[�޺O����/g�nj������(��#�K|���ѹ3��l��~��}�sv���FK|'����1;cn��H_a��D>�h����λQ.)�{ ���YeX�鉀�餽ܮ9�?����8�,/? ���ρn���h:���C!���(��#�������q�}X<G�ZGtq\���Jj���$=�~�ў��O6^Y|Qn��vS�;�߸?m��K����޶�\It�O���w�'��p/��gjw��j����n&��ڵS����'N�k�|�o��o��z7?�u�i�Ԧ�U�������������C֭L�u�)��m2�o���a�u�ƛ��Q�z���f������6j���<��w�o�����B�?�K�<�}�G9Ӷ�EVq�~'(�����̟|�Qv�8�!:���?��j��e��&��_��7ˏ)z_'�O�Xi���R�������t���6�g+�����8"��`q�8N��6>��k˗���yef�������2�n)�����	��ɞ�?tX|����/^����G�e^z�;y(��
��v������5�[d�o��������ٸd����W*���:���L��e�E�管�Y�[��3��)�3��?��x�>{b��Y��K�,{?ߋ��~l!���G�����q��~C�_D��e��5�3�{.���3{ש��?��~���?����QQ�"�~V}�{�,�9���1;O�}�#2���~-Η����nYőQ9���c���	���~B9}~ͫ�����x\2�G?_U����[�33;����U��Ԯ��ϓ������n��cϟ�o��'q|*�{dxKñ�l|Db=�o�Y����S=�Vyg�%�_��qvi�=_���������r��K�3jҳyhv&���ײUG�=���˖Z�s���اȾ�1���YY���7���ϓ�c���f�V�W�����6F�������hF������
��_���o�?c� ^w4mJO ��0�ܡ݉��7|��d��}�ŵ�v�).��d=3�z��m�w샖�b�����\#_��e}�����.io~�E�9_.{1�uo����3�?��'Vޏ��|�s�u����[���?m����2���C���q�t]�%��9뫬>�2����g*M�����l߭[O#z��q��1��u�)"��P~����W���~r[��l?��ɍ�+����E6���]��Z�y���w��9�o����st���1|��G7+�E��5/���~���S<�y�����f)�a�]���{L�I�y:Ɓ����N}R�]/��n��fmf�|���g�!�'�������Z�?�ү����>Y�'�OM>���=#��fq�]��&�o<�(���{y�f������o����ߐn��o���u��Ӳ��W�3�$��=�?*�[��.����;f92����y�����lً��'����J��y�4�I<ӭ�l'�����?����2KG$ƣ�}C�9ψn��?���Aph\O��ѿ�q����G��7�����C��?^WI<���'
���h������>t�>G�C���r3<aѩ�Y�Ζ*} ���s2��� L�os�}K�M��=���L���9L���o���zm��nԽ��=�ڿ6���J;%m���:F��u��M�'��`���������+� �ǔ�۬�G�3�s7�7��0G-~{�Se�R�X�e��ָR�������ۥ�/�����7��Hﭣc���bN!��䢗��yPL��mR{��5�q����G�2��^��M�}(ѹ�k㾛�s[����kM��~��[�-f�祔�b���o�<E�� x�������=�'��Sz&�s���Z��J���9	=+7jW��ϯ��c]$��z����V���C���3�ߴ��|/2���W���o��z�1�2�'��F�N�/����:��S��"����~���.	=��d)���c�x�?0��Y�y�j���]����׻#@k9'��t���36�4���Ǭ�>��0uo���7���G��	������kdxQ]/�=�O��J`=���*]}'�A~M�c�����#���G;0���<��5�GR�G�|O'��c�������^�Z�q��A�o�w�����h���y}6{��;���a~��"c;���7��+�Ӑ��v����2���ZG�G�٥V6�L���os�0j�o�?��u���ei�~۫��=&�}��ox��΋�ه�?�Gԟ�O%>���k����n&/�zv^�@��l]�����u!�o���0�� ~EV���ٺ���2�oz�W�˺�xg��
��('X�̮���֏:^ѽ�M�g��Aq�H��g�������>����O�6�A��eg���#�Ǻ�;Dz���K�����_S����&ۗe���}��/��2?�H�_��\�ue����׈,^�o����%�M��^]�߷;��9���#?Q�o������6�F�M�Ga���~��T�x�g��~c��<f嶎����&�������2����zN��`�ټT����o��H��
�{[v�g6����}�K[�A�՟q��d-{��זG<�p&��ҡ����@�rq9�g܈�7?ۓ6�Z�Cfg�>�p/S������wUˋ�7lW������(�Lɯ�9�cG%����s;�?[/":�G�"�%*��4�3�[g�F�l^�8ۧ?�>k��~$[װ"�yf�Xx�K�?+���,w�����L�{^Sq�2;D��NY��zDr��е���Y̹����?��qc.#y9���O,���(�շ���s�������������}jC�u\�Z�xN�|�v�=�;�1Q���{��_*�8~7���{�u�Qb?n���g~B���.�y�����w�x�̮�deM��h��]��q|`���ҏ3�S�G�� f?g84ƛ��O�����6��z��Q���ƣ��b(NB�t�%�W�V|���ˀ����i��3]�64��KdK���1��Grgm��|�4����>fx9�?����[˟����1��'�������E�ӏ�o+�5&�C������8�H^؎='�g�1!�+��"w��\<_S�����o]q��	���
t��u��>���~�������>�1��T��-��4�%��e<�~�f?#����\߃��k�O�|4f��&�@|�M�˟S=?���n�����d?��g��[���~�>_%c�df��>+�Ň���On���<�Xk�Z���s��\O���u�#܅}�t^��\>;ύ����ؖ��~�������keW�����_���oŽ��.��S��Da���>�虽��U���߻� ���oG�S��b��6�ϣ~�JY�������%k�a�ry~Z���c���[������*]�[x���w�=��0ړ^K��m��u���yD�����y5/��G���G��k>�W�~�z&�ၿ'r�u"g�[���N�"?��Yj��Y���c���;$�{#��˽Tb���=5߲�f�<��5��a�o��`�����޲= @��������OVϖX���ϥ��h�Zb���gj������\>�Q~��������1��_�Jڋ�c�lGevB��.�ʆꩿ,��O����_�ײ������N����q�+:}㮤]X���s�)���`����%�џ�W�A���Wu����m�_�KF�������$?��6��ɸ?-mJ,_"�9E����czG�M�u�Pޭ��x _]��N�v��03����M�/���v�������>���xb�r�Qy��|��d8|�Ϩ�u!�i���Ӿ���`��1����~乌��~��[xmM��<�3���[�g��u��s��/��?��w�N�EY=-eq&��b��~Z=���ھ�|Db}��[�?�����=�?N�q�L�h�Pާ�W\{O��2~�R�ߟ�_�oh�|{��c�ϙ�g���z �D�~6����t��]X!�S�Z�*��m����\�grd���Q}��|^���	:�s���n�_�Hx�厚W������0n��c����R"?a빃�L��wS�=���ůc?3��%��I}���:#�u
��~+˻����T���U^��9����;|�����G��~P9�q��U[���Zf�G5C�'d��+��I���<_������~��X���H?Yi�&>&����y��s��o��R���eͧ�/��������g	��}��-�gN%��^��8��@t���/�k߇S?�^��q�%>6�L���8�f����t{���d�]�	���fXw	�,_v~������⠦�+���t�tG�?ڿp��O;w���(S�˶��e
}w�?�g�O�k�&+���!�=��ۯ
��~�1��u�y�������l\Lo����fqKlnG����&��}�g\��a;��x>��W�M�l�+�s�^K�.��.:t�����ŵ�w$������:��~�Z��j�^�
Y��F��M�����
���Jמ��y�%������r����ye��A��d��������%�o#]:�L.�7��M��˧�i���T��9�ڕh�������G�JY?�?*Z/l������w����ڗzn��@������
C������Jg�������u��3����~����kx.cv*�=�����f}���%ާ�X��Ɩ�.YŖg��za�M�7㓽G��;߃0|,㽱.X�߮<�M�y8�yx�'jo����3���5�ͺ��&���6��E�y�i��G������-��dܟf�fqy��qe{�N-�Yl'��Ϫ�M�ߺq���#q|���>�i�}x__�=�ZY��V}�Yw"��
�c�������`v��+�"~�ՙ��_?�ߤ���	:���!�5|p�l]{�����g��[������yI����]�~k�5�{��:���$����o�5�����5��zu����cB�y��<�{(0���s�l�^G|2��7�
��[�C��F>ܧS����������gq��sR���@� ?ӳ�S'���9�L?�R�]B7�a�M�>�^��'���+^��-6ٟ��'����&���X�p]��E;�o���V� �}Ǽ���E��ȯ�?|���V��|FqY��	�=ˏ�<U��L�g~��O��ȏ|��E(F���D���?f�Z�]���ہ���~�(�;�R�x��ǰ�\�O�����:�����}�h���Zb}��G��ջK����s�'��������ݟ��J?!9^+�c����O�J7�����y��O����'�>�����JW���/Vy��=;�H�x���z_^��3��^���yxRb��>�����t���w���o�ؕ�;d����U{壅��Y�xd��[����]-�0�Z�en���$��?�ʽF���!z��A��~y~"��@?&��sE���������Z��i]P�����}��W*�=��s�\�~������u�����hQ�-�e��s�s��A��0����%��T:���m|�|���Yuk��^�~e�������(��؟c���Ք��U� -�d�����f������݇2^�n��^J�T�Mc����j�"��������e�on��D����U�<Y?������2�����f�b��^�������"��ۧ�g=È�*����B۫�g�-��c������Z�S�-kW�'˟�g;����Ww�jL"�-�'��`)×f�'�G������Ѻ��#�翍����;w���\3"���$���߬>�S}ʾ{ϿyR���)�}�X�Ӳ����X�?�?�h��v���p�CL�5�o��l���\t���.������g�+҇�:>�����o��۴�OŇ�KVv��>d�n�zY�fE�E�m-�y�������[��l�׼g����o8�����IǏ�s�S��+��Fߪϛ2�?����e�`+>
i-�J���=�I���u�e�оz��{ә�F{��	����:f*�O������3;�R�Gۖ����A�������T���<���5�H��ͫl�]�"Z�2?jv��E�f�A9��OE�S������<3��_�D8�sP=?����H�9
�6{KB�;���?˅�\�9�!D=��/��Aἲ��-D��X������:<���啶��?:�֤��S@?S�/~�>}�~F�O������:��LY�,���t����||��k��_ �{I�Z��8?#�M�^��D?��|���r�=�����W������x#��f���I��b�y��)���{OQ|Nn��7Ø>������};��j�w�y��S��q�3�%�����8�(�h]�{L�K��ѳ�������fN����7����9� ����܃�Gc���j��惎-��V=���۽�2_f���{g�?���Չ�G��}h6p�mqs��Z�s��%�C�N,����?��+e/}���s�f��彦|��K��p^������2��Ŕ]���=�Ε��x��d{���nּ:�n:���#��s�[Vk������C�!ֶȾb=`��h�k_��#�����g����m�x��P&���q� {1g�������]�S��0��7�O|M�S����8��O��&�����Ҷe���=D;G�5�?���/�3�U�S�~��&��3⾘���]?���<��޾O���R%���X���fI�G���De�� �:��u������-�g��T�Bo�6�T���O�F`�S��gԇ�L�[��	�2y7^�FW�8�=���s$��ۗ!=�m���㉽�~���&�Fz#�ϭ�m���2���}����Klwe���3�C����?P���-����پL�zr�W�zk�������>G�j/���D����Ke'p�O�������$Y?L�5��������>�>���� ��E���t>�'󋮫'�����z���/�?�;�}�=2�?��K�;�va�w���e������=�{�X�WV���i��+=�?�no�o�'�na������'��W�o����|�>O�Cl+�m^e���5�����A�,~Bvn�z Ç[��O��pk���xѶ�s}p�G��ռ/�������E����2S���?�<����S��C�ϵ�����=��-�+Ϫt���TO��2~o�D,�ڼ	�l�0unh�1=�7z�ң�i��F�|(/�g8J|,�$�7����F���q8*�?r��;de�]����L>ٺ���?y,�#D��'���-.$�u�7Y�8^w2\���Rʏ���9��Im�3@���ݯa{��e�_e�+��3�ɺsƖ��q�Z����D>&ܟ�����4ǧ4���l�~K�*������7Y?@�^g��ګ�P���e����/�
���aV?ѯ�����G�%�?���O�/�� � �Gz5�qZ�j�b��l܍����`2��f?U��.V>1n�%ܲ'�i����~K��7T���B���V �7�79�8K�XO�o�oj|R�sk�'����g��Ke_f��:X�T�	��>}�y���㜣����Ӳ�;>�ʽ��i��~���%�����ʝڏ�����x$�_R�Ω�}���e�ް�]�4���d�Z����.���"}qf��F�7�t|oET������P������=��������.�+�2�����!ߧ�t��>�O�������?~����%K�_��x�evHƟ�[t���e���?@�V��Ж�K����)S��=������󨞭����-e���~��������%��3�g��u�"]u��du��m@�8��,+���|��X�����O���]��3�������`/��իߺu���a}2<ITO�O���!ң�8����zV��U�um)�������f8F���5���^U�NƸ�)?v/T��H�[]��=�ӟ�|i����E&��yt�2=��?�S��o�>���՛��8�qD[$*���i���ϫ�d���ߦڋt���+�W�j����zZ�پż\�j?��O�=pic~՛�տ������O�U��s�_e�>�+���L�����-2և&'��s5E�׭������Y�����t<�@�}rć�)e��S8�.Z�#��%�w���D�9P�z��2�Ge�[:�+��ߔ�<�����sS����ίV�,?)χ���w�J�򕬿��d)��eh����{���*S�!���1�́~u���ը��7F/��޻�,��qA��Q���n���}�mE?	�cXO孱�to�簘p��nн��k_������>�zs}���8��7��K�+�Z��K�k=Q�G9B{8��x�=)�}��_ĵ����L�5�KF��]�Gt��b�M��k_񊑼s���>�L*~�����=;����̎���d1���|�K���sӷ�&������i��D��2��>W�����z����2>����x�X�9~�!������=��ׄ�5kov^�z���������s�uq�����k��\�������踿��s��[<]�N���F��N�x�Zp���+�ʖ�?`����R?�u!_��'���x~Z��[�n�,}wG���d��tT<��@?S�ܿ՟���HW���E�^�kerar�|p]S'j9s���Lϥ��f�G�W�/����g���u|0���N�x}�~@=c�U�_�_wҢ?/��x��������-��fx�d��qf�%n����w-�ͬ���'zv�b��~0^l�X}���x\����|�����x���t�s�>d�ͷI�\�S:�T^�B�|`�[fw�����z��y���}+{�R�ޡ<Z}���!�po�U���d��wI�[��s"��ѽ��T�);˝�Q�q��Ż�x�Q�p���t,w��Í�bX�lߊ��u���_X���?�ڥ�.�o��ۊ�A;-�������>i/�kr��O��ƹ5�ư�>�+�����l��&ȟ���N����i2�?��:���4]GU~1�nV�/��=�bnD��̞�I���=���w���tnf���t>/@;��c�T�����:^�R��}ٛo�{���.Z�zt�i�����v.�-�����}|6���u��-^5�g���l:�>OV����b~%�C�􃥉y����d��-��A~�O�E���>�+��q����$[���u�W��e}����1��)2^צ��օú��.����w���d܈�7�}+K<O4ߗ�ʎ�M�gzە��~�6\*�{��Ƿ�ߥ:�ɵ���<.Z�_=I��e��$�K>X�g�M�7F�}�<�!�%�1>��R����g�fğ�kߝ'����%Z������T���I���xq=u-xz����c%�?�>t�{�����������ڮ9���uG;�D��I����r3��vE��}��ߠ���T��r�Ѐ�����^����G��k=؞�{+(�g+m.��\n��fLw��Ν������͆���h�h=��?*+LV��3<����Ӏޗ��aT���q�Cͫ2��+�a���7�
���8ff�\"~��g$_/�>�����b?�������=Gx][_-�y.��T�}��+G�W���˘����[˾lv3�=qK�v�@�H�?�uѹ�/��4�~̽�Nx�ʒa������C�<�/�[ڼ3�u�?{D�:h���o�g�G� �7}�Hj/��c=�nv�92�W��2��|U����}�쿕?}Ei�^,9/ŵ����+��aC�������oW��3;����K���������/�������-�]�qZ�����~�ΧsႬ�FZ����yG�ǳ}����T����ُ��o�dl/�{���7������k��d���MGk>�W�Lu�A�Y�Ϫ�Q���P�C�MV}����"��2�~�){,;���|_�X���|�Cr��b���u��8Y��_�D���⯳~S>��gt����Hi}>K��y�w��}2z_����[yY|^���l�l�w��������_��n�gv�ʢvٹ�W�shշS�֌�A�V�Ժc��&��m�s����<t���56�<��s�ټ�u����@j�j��U>پ5;�8U�R�d�Ǆ���G3촌�q�/RL�q�+D{��B��御T��e�ޥȟ�m�D���2�_`�T���>��p�{���W�w��G���p�#��&Q{M���o��pPz�a�����ɐ�Ӂ���e�'��sV��o��Fv����WS��/�{��/�� ?��Q�K��0�z��\���].m���R��c��Y��q�Y��>}�wT�m���R��?���Ogܿ��<����D��"Gw�Jn]Sv?��ۋ�7o�s2z��Q!���V>��}��#Տ��u����S��:��\.cy����	>�����]2���U���"���۝N/��J��LcT��R�+���!>3i�����O�x�bz��0���3�vV�w�^�\���y��޿�;Wc4Dv��J�X~�U�sϙ����K~�|�]ȿ.~��7^ٹ3����D���ev���;�Y,�g����;Et������6��ሲ}˗�W�ߒ�?ꓬ����U_k�= �o��r�����4��]�RnFW���^}�� ��_�W���'��������O����z���������/2^<��oo�3>��f�:�yU���q���=�Ѽe�ڠ�L���ɿ�ռ��<��5'dA��uZ�K�������jl��jӛ�W���`��U_�e/.Yp���8'��vB&GY|�l�0����������C�m|ޚ巔��~���'e��B���$��|�m��z������+�X��J��f��KV�Ï�����e�Q���_��? ���l��8��܀�uD��ů{0��u<*���Xm����3�F�9t�i��#|�Y���l�f���G=��B������tY}2ܸ���fܛ�����~B�����2�k��i�˵�H��C���������)�G���yk���@ȋ�&�;]\��*yf/����><�2�����ZF�'�'���X��_�q�R�uR�<������^i��r�ߎ�O���c��'ד��՝�k}8�oq���5��Bt�N�G�#��7�����h޲�:�v��e_W�]d�.����ߌ�{��}��u8��J�<���g�/Yy"z���������;��x|����޺��Z��|X�� �������9���Oq����)b<����������\V6ﻳ�L�#8�w�g�/�is��Ì�n������������O�J7|}C=�M�����U�)��a�����q���S���*�����l8��,�ir��Ym����˧���&+_���_�ο�^���`��h��$m�
�G�֓�"}N�������>�i�}_.�Ӳu<�!�����Ѻ`8�)�B�M��������vo������#�q�粒u�1�)����t=B�����5�s����u�3��^Y�ˁ�P���c^-c�7��>�uV��Z��A}2�Ჹ><-�G��]�A��:=�t�����|���?J���Y�@�g��DxN�X/���Z?�+�?<��\�36�'%�����QQ�,C}~����ں� �g;W�r�φ:k�߲vY�<�2\��+�������$?����N���f��˟�3ҳ�ۂ������u��X�����[p���nv��ʔa ��7g_Y��҆�Y=u����&�g�|V�}�@?!�1xX-"���C"��L����k�����x��q�e?��뭲�}���ه�J��G����]��wh^�+��lO����}�+��HOf�mC��q\�m����L�ËZ�ګ_"��0�� �c(G(�	���eu���;��n��?��l��r�sd�w|�򛞽��6ޙ?��Zc&�.T���A=Y�Y�0N�b��O���վ���C��ng�����a�6~��y?�q23{�Y+/G�}���㛭��x�0.�� ?���St_�!�^���g��c6������#.�Ϫ�0>df���U&�3]��W��D��k��+���8Y܌����0�걖���t:��)~�g���x���}��5���xd);O��#\��j��g�1�R�=#��[��c��s�c@~�){1�����q��s������y}V;�;��ybz ;���N���>���)�;���������of�ufWp�B�׷�s�G��j��d?�{��CT��M�i�Y��6�,/z���l}��g���?jS������е<����qz-~-˻��g��u��r�����	<^ǁ���7>�?��;�p?X~��cJ�~����T��{��~����h_
�����9���:+q�"���w����/���|}g�D}�Y��8���s������l�^+��m�����Ez6O��y��vy�ʽm�w�%�ױ�عcf<(�����u9�W<�&��[����g|��߻���h�r_��	����MOO���w���]�N�É����Q��?Ю3{�a����?�tR�V<�%���|����d���~P=vqm����ۣ>�%������}�?��Py��k�����O�umyo��C�_�xΉ��}�f)�=&�V�/�#�s�����c����8��A���v��S�\@tLS�>K��گp�{V�:�^�{w��&|Z�=��h�Nq|ō$������P�_@����xCC�m�t�\���5���Gy	�OԼ:?O7����M_e�y�������������c�_� �#�>�F����Z�$���bNvN��kC�S��b�c��w��Q1^S�\ N�b��^D������V���)��u���<�^�~��}?�3\��7�g]�"=p��I��������#;'�vi_++ym�����#���O:�Q��e5���ʏ���f��+���Ƌ�L/����'��*�d�m!����}p3��ĿM��<)W�y4�|~jr��fq�.�8>��c�7��@�(���Wdu�O�	�?���i�Kڞ'�g<'����*j��{�X�e���.m�o��c<��f�~�&�5?�q�s�'��2yA��m<������9ٺ�����J�9�7���z�[�g"�xފ�'��?,_���H��/��j�2?ɺ���\�Y�T���8)��#Z���?��֥��g��d<^O��[�{��#,�9��G��BtK<oߠ���W�]��]��Z4��=���\L<���W(��Ǭ�R���>�P����j�t��I�XıG����}[溆�/���I�β�$��>��ǯ��~.�#2��ϯ�������?������j}��޿��GS[���.��L�5ܧ�e���	������)���J��������A~��#�o<���{�����gʎR�}y^�Y��ò�kւ�ڀ�C��!����kdkS}C�Ӑ�
(;;����{�-������{+]�!��2��^��=��]䷱��c�3�������0�	��Z&��Z������ �~�l~ںr��[�q���,��k�����_���'� �9ڜ虞��Y�9��;e���N�yxn;�{a=���3��ߔ�|0�o��Ժ�4�?z��m�c�P}f��ug
�s��z���~�l��_��V���g��yPO�oi�����H����J�7�<{G���=�נ��t+�ϣ�������@?Q�K|�%��q�d��I�籀����\�|h�������Ԡ�·糕����������yk��N]�7�KV�F�� ��\ۻ�h�s�XK<O0?�[ܿ��d���x�gx�YR�.���f�eX���,��������{@RO�P��P�WP}P�_J�LNm\�C��e��.�C��74�|C���k!�]����� ���z�Y[��$ϓ�����ߏ�I?*����P>��|��Z��
���	���4	����g��]ъ�B�H��>����˟'c=���'e��>��JSϖ��O�#Ɖ���+��D��y��r?`�Ƶ�#+_�x_Y���1L.���V�[��S��[����Y����[~�؀O����)MQ������|����Gz��?S�q�c�"?g��˻틯���]�ϣz�������q@?������v���S��Z�zl�߄������/��xV���4�Wfϭ����o��5��������F�1ғ$_�?�|�]�w_I�uPꇍb��Xt��g���	�[�?;#+{�<����m�Txc!��5��8�P��{�.�<^S�W%ɏt�t|���k���z��v���ٹF2^{����{��7�jo���}��HN����끨�'���Ǹ!�	���S��%�O"�,���oZ�5�)ϫ���~P�;��d�����LGr�Z/�7̯�~�=ԗ=���&�c��8d\����"~\�<��TK��e��0e�6����H����~����X�y�q�Z����Q���2VGT�[a�� ���~��ǅ�\ß��zڸ�e�>\k�#d���QV{8�K?t�}}TVs.:��q��+�g�R�����a�e<0�[�/�����Y�S����f��-�#�/��:�'���s�t����k7_�bM~B�����ƅ�c���/��bQ�����׵��d��ҵ�?�uV:�歕mz�ʧ�"����o�묝S(�@7�����Q�p��g2���곞!��c+�C܇>q�9S�;<_��fo�e�v�����������<W�:�����}�!�{*{�2�7���xѩ�o6o��H�>��x~b=��Y�Y����]|�E]_��dV6����6��%�۹����=��W�i/ӳ�֏�K��M0�|��e<�����g�	e�3����՛�"���{�Q�:7��������fv�0�۸�N|��7���}d�Mh/�s7h���u���o�׋)�'���0e�$���o����wK~�L��	�-����o��Rv_,�O�^�:���r��>�O��{ُs{X��x��A~�'7U�T�.ί~�\\E��Y۝��g��oO�*M������_�!���`{1��!���)��g;�8Jt�\	߳^j������M�]�c:^z֍�)Xả������0Z/"z��4�|9�w����{)�+X�g���5�G��뷳�v���3���7�w�8G����ML���vJ��4��x�����4���#�l]�2#���]ﳨ~�&˯̓�����x�׵�zf���W&�s�O�����Ӳz���u+�Of�>��I�>�:t�vF��-�h���VBv�g�ﳲz���^ �^��ږx������f�7������_��9�fUm겿�E�����߲�����xiͧ<z��WV�T���ղ�����-?D��XٺO{h�i�G���9�g]��vP���5�O��7����bW��ɷ��~?ȟ�{���xv�5���ޟ�)���<Y�7�~�>o�'��=���w���7ʞpC����\8����Ef�����-@�}֕r�}D��Ь>Y\z^ߧ�\�E�y�M��O��Mח��0��x}�D�c|/%��c���B~�73��w��U���/|��Ժ�q� /�Qʛ)���J񈷱q���ZG�ATq_����x\�ZVsJ�wď���Ԋۑz��.�6�Hʝ��>�����s�����#�������S|�;���q_$+<�@~�:]�>(+��a�����m(ϻo�u�XH����]�x>����m�0<&�aQvn;U�W�{��!�1��)�_�G���E��l�M�[g��[d�����h���s��X�� >���C��g���CA}���3� ��evL_��4�Ǯr�����ϩ������s����9Y{�o�d~���)v���d5&-�q���������5�o��-��T}x|�U�U�����M�xJvǫ���]w�sUοY�?�����@���F�O���濎g��ȳ����'����Z�(�dtbw#��1�uo�����@Vg0*�x/y!����:P�[��Kۺ��s���%2>*{�ktsy|1�ͮU;6:���i��oHG|�;����z,��p��|��������/-E_
�m�8M��8�x�h�v�>������֠߬�0?7����H|�*���ȿg��^s��O��G$�Z�m�wϗ��2�Ǿ��#��+�0���g&�����?f�h�(��P�"�3�_�k�6��S��v���w��1��Ymz�c��x�*��n�p#���cD�y�Uw�OE�.���2������2N���"=G�7�=�|�����=����G��_./�"��g�O��e��֩,?�K1�j�����@���X����χ��K��}���m�=bM�#=�x<�����'�����������?Jӹ2>/����6���!��X7��y���[�@tۏq| L��b}n,�:��*~*���	�g�>I�S���̿��i�a�T�<�-?�����SeQב�}���b��>����g�����?��a���6�����|@�m��ۨ>6NٹC��f�Y�e�rm�\���	��%��m\���e�/�/8++�Ku��>�Xoh�0����.���	@G�Gt+ۧp?�}X�g�^ij'>G���6�`-�<Z��Z}#���2��8�+�?q�c��rvx����BV�ݝ*����5ʝm���i��l̩��X��~!�wl��|�����o�>�~">6���vo���q��W�x~r�K,���~P�y_-��~���6���~���B�l�iz�0|�:�}����y�zb}>M�����+���v��m�x����<&c?��<++������Z�O����D\Pv���W���xI��(����S��l������/��p�>}^�#����C"�9�.<��n4�0�A��W�꤬읻���8Z��oz�H�V��i����hYz��(Yݩ���?�{���r��˽N����5�k%����m��εYџ�7���!�;Y醧|��p�m���Ŏ�5���t����s���4�����U����d��+�O����f�������X�Q|i���G�3��d���������^�֣);��[j=�9����/��8j���_B?����Aֻ��,_��t~��&��>�g 홨���<�t�G��ߖ.=t��h�(n�����~�n(��#����΢"��z�i��ϕX?�>��U[��Rf7b~��[�{���f[�2?I�o��g�{�c�_:�A=�~L����X�;�۔���~CBT^O�ޅ���V�)=����/��"�Gt�Z��x�6����%������M��~"�g�_�'(A��	���X�����TL��˞�f���̿tk��lY�� }^��8D�ϑ-�`�[�~���<O2��	���m��Ɩ���Kd'`Jj<�_�=��C�2�D�<^����`*�hȟ�k�|*����1�t��k���ϓQ��{�����?��/�m/�<�!�;��f��{ٔ�9���Sm�?h������3m�r��{4>?���(��w�x:wH�������ǑSl�������n���8?��R�g6�G:�'�y��-��v�=�޶��9N�'4:�dl\7d��|�9���K�zfz8kW+]׳w��;E�poftۓ�vM�+�3�V;"����g^��?��ꗺ[�8r���O ���K$�;��g�)���Ѻ���>����҆�� ��ȇ��K�7����*W���f�iz���}��T?�Ϫ�#&��m�Y���<"�g��_���o�~�\Bt���x���|~����+��w?��gk~���/�G���ˋ����[�,E���u0ñc�k��}ٟv���<��c[�z�wS�֒�wt�bu���0��l_���|�n����o������,�V�<iWV�K��G����R�ϕ,�5}���s�g�O�^�����������UVwq0.����א�S���e_�y��u��ڎG5�q��Kv�]m�k+|O�$�-e���7�v򱄞����W���'ٹ��^�O>`{���+��4\��Z:�}����pz����h/��㈸�S?�"+�F�:�k��A���~��5���+]�����`�y��ʢ�(���;�	����3N��W�� �u�jW�9����~�躯��<�w��f����W�x�u݊�L�p]6{��k�t#�_�'����R�j_���q���4ѳ��x�\(�{�{�nv5ˣ����)=�n/�3D>=_���ّ�w��-�y���	�'�Y]�� :�ۣz�����F'c��e���Ju�������<.6��x�0;�@��>�]�z���4>铠ޘ��,��:�eV���/��JS������I4�׭S��vN�ϗ�J�
�+���.����J�����R���y�v��������q���N�6T����������n�o�ϲ���~�>{Тr���[=��@�{�ϗ�w�p�l.D�=Ⱥlrܲ<��޷���]i�{��5�F\�Lu�o������u��s&G�N]&�10Z�<'��F���K�(o�|����d[����l|�ߎ��u���ʜ<��{7�웃������"{/��}���u��Sd�e�d=f1t3|o�'�ۉ�Q��s����������A�d����G��-�����{`3�{�L�<��U޵�?zor�#z�Gj9���k�믶���3���?]�����r3�?�M�n㧶 ����l�G�2�3�ǐ��
��o]�.�����5���o�s�l>[��	���cV�4{�������:Y��7`�ؾ��ߟ�����[e�MXW����"�փl]�u�ΙN�X?�u�{a��c����ߣT.ƝC��ޣs���>?��p߱~��d�����3�W�;++���I<�x�������G��Ԣ絟�OV�,��|�m�W�H�oy|��x,����ֹ��a�s���@��~_V:�ր�a��O#�`	�&���|6���^L���S�K|�*��� k�	�k������d<.�*���G1��=o�����ֽ_���L�	�D�S�|f���\�~�w�
�g�(��~k�Se�Y��O��6<����վ����읫o�����:�!,�خ�F���/�}�����a��h�x;��P�ras����W�%���LOF�u�C��".�_���[�!"�i���F����"�|���3<�}7eg�@�]��,�xD�^�y|3{2�c�sC�q�z����e��O?�=E��Q��J�~r�����e�;��R���}L�uA����Nv��}�����	�>Q�ސ��ҧگ(�-~�g������D������q@��55����y���!dv{��^ 4��>�<����Pϕ����3���ǈn)��&�l�g�l�7��ג?��M�kk���#�*�A�+���[V6��l����%+}��*w��D�)��5�ڏY<a���1�ޔߕ�.���:Y�k�����[L�r���觠�6��x�����*]�R��Np�z���<Գ�{�r��?eON�-�c����R���|�p�؟hcE��h>pBKl��j�����L�Q=)^����z��)�.�ݺ�8(Ŝ�ٕ��S��^���պ��n�[�š��<ߌ�S�?����!���9��e"=�b�~�������}��s���r�^mݧ<X�	�����_R��@;�C��Ԫ.�c�Aͯ���D㝪�v������\��lj��xjs-:����iY�uL�'�p���\��tJ�dr�)�8��o�?u]�߲g�΢��G%��l���St< ]�I�ߡc|���e]���a��Y�?�=;�b?�T<�wqP���Q������R�Oߟ�~�{�P~�nl��c~��_k�ᬽ�T�������T�� .� �v�� =��0�����dv��E�^�Ƌ�s�l缜���'q�q�Ε�;��l��/�����܌�=�-�/��!���v���;O�B�5;�z�o�f���}������nﺸ��6���'�EV�a����O�߫���ď��x������?P��粺�'�"��j�f���m!��/����]�wz���A�\~�aY�5_���-��+}�����ߏ�0�������YٹX��4�b���~�����7��1���2�{6o��ٖx�;$�غe��=�.e����e������v:v ��$�'���-���{���M�g�Ӗ���&��	��l\0Nrw�yK���-��2?�������2�Ad,/�Vڷ���W�X�V:뙹�����?#�\����q��~�x���;ŏ�Q�	�;����NV�T�l^i|��Zt/��sA����J��гsjK<�����dl��:~������Wَ�da�-�����~��CDb��z;�_i,�-�7��~_��,.(�۬]*_O���C����R��r�|,q?��zDb{)�wd�/�Wd����Y߿т�}E!�]�����e�X�7o
����տ���7�������}����2ޯY�d�.���й���@7��ש��_6�.������8���)�2��뙝��ofҶ����K��o��m��ҿK���|8�S��87�~����@L�z�����K�ù���p�Q��U��h�O�.ӧ7&|l���l�ٞ9Vy?T6���Q��L�dx�VyAz����'R{�s�L��<y���6�����sRVs]�;��Rv�հ���� ?�k�\�d����s��o�g=�ޏv���O���3�k�ׇ>������/�G�r��J�}=��e_Fq\Я���O��i~�J.-�bK���r������u8
���ݶ!����f��ȏv���MTm��C�����=r�xM�zt4�P=��=�;+�s�5����8�����T�>�POۇp�l��{�q������Z'��Z� �}�,^������!�+�@�]��[�-e,w6o�8`V�?�W��#�+��w�I��}��g�_�L�������3@7�=&c\ڟ-��Wi)�W�v��4�9����tϧ2��Ij/e�20dWD�\����u.c���y�'��yN����}��
������u�Op>\<���9��⴨����_��������^'�{�V����q#�~��Z��*��yl���m�c�q�Mo_I|,�Iˑ����ʗw\��Yw�M����QW�����f���g�>�_��x<��c�}�)��e���7��k���g�{�o�&�6���Z���g�N�cٺ���;����*�o�׽'(�kw��g�z^���}\}�xV�_�rMN[q&��D>�}�\kTn�W���"�r7�N�w���Yt��4�<G=i�@��}ǛeͷV?��_}�s�ש,>6��]f���3�?�ǆ�������~�rͮ�q�u���:�F��>���y�iq\�\U�-�&zkP�s�>�����T:ߟ2����E~��\f�}�B�~��d�� ���,�\g�������}M!?#(��:��v��m��~h��������qe�r��4o,7���]#z6^������[/��Я��i�������wj�t]~b����|������(���35�D���e_F8�̿'D��N���р���Ѻ��v5��6.&>�e8.����8�����ΐ����Sc��zs���A쇙��+��۽�����d�������=����[�q��>����{Y������l�[����a��M�c��_��5��+���5�3\�b����.�����hY���d���8�:�ٓ���9����~��#�� ��������������.�'���u�-��kl<�~�+���y���t�������k&Z���[=i�7>���*�Y������Ke� q���)�i}��<���4{����Y�?3�Gsq����|�k�R��?)+<�T=��� Gdߞ�r�7s���揭Y��8��Q?�ްy���pM� �cmc�b�����ݫ�t�<a��cz�%�k�����Ap8�e5�g%��c80�%�M��p��d�kgo
�D��>��������������4�/��>D?0���^�g�]�6/�a~���wI�����C�cc|
�o�彚�[�k;6�nzR�#������� ���[׊'�~�|��j-Թ����X�{��\G�DvB�Wѻ'e|k)���_%�a��>�|��n������-ӫ�~��):��}j�����U5/�7�g��#>�ε����s�~��}�ف��x^6���~F>��d7n���]�Zs6Zp܆��9�޴��-�=���ё�C��T��m�EG�F����>$*���7�g�^K��x|Uߝ��\�%�!|v}V,�ۨ]�w\�~f�?vNn��N���M|�<T���������/8�����ډ�ѻ�O���iQ~����5SzO��E\ c���3��Z���Q��WB{�}u��J1�~�G������Z�=�&/�������^YaUm~^Z���R�q�~�'��;0�C�O��-Ok�6&�ެ����Gdv�Ճ�}|gy|��|̈�ȏ|l�=&��/�z�"���ѱ���T{-�(�ov������k=1�@�!.�S�K�jd�Fv��kğ��\Dy/r=Ӿ��HO�ʞ��;V���6hov_����d%s'���z��g~��uV��!Yټ��ʳ�[�'�U���r��yF��]A?�O[�/����f��~�����]�Z��Kl�����_��ߥiNt��(��3_++B;�Z���U~�㠾�g�O�7g�Ηx_#��4a����s$�O�ٙ�������P�cB����X:�'�yk	�G�2O�8��Յ�c�|�+��L��ӷ�."��~��;Ob}�uA�o��X]{���C�퉀�U����w��������R�O�r���1ęo�u���ҍO��vJp��/og6�.�������r��-�aK���������n�����1��~�n�,+y�SV1Nﯽq�>?H��������}4��x.�t���pgo�=�t\�2<FT�u��H.�L�3����,��~����A�������g�_g�n�����fq�n�
�螅�W��볮8����t|o�p=���
�~*;�P>T��_�=,�,�;��3<��<D?UT���<Q=�~|^G��qfl]���3���&�S���q9Q��J|^`��M�Kƽ���z�������Y���,��L�Ⱦc9�3_���F|f���_=)m��S��v���;��f?/�����+ڕ���ݬ����ۍ�����BG5�Sො���{��/|�w]}�>Ƹ��_'e������wǶ��[�[�?��c}b�~L�qn�<��;�Ǒ�
ۿt}��_֓'e�^o����>U�눮�f�U���k��Շq�jӽNV������Թ��#�ǁ���3-�G{��l�T7�\dz��`��K[tO�)���k�1�w�'��uvr�g����p���8��߶���#>�ϳ��>����tm��R}���o������8��e��{�^��%��xN��6���J��f���O3?��V�=�[��ox�q)�U�Fѩ��پ���a�G�d;Ǿc�d����-M�[���;��d�M�3S�ʪ~~�1_W�W�n)[�y^�9KDg��3����W��ғ'��"=��������?���������%_��;�ٻ/�����k?d�PK�۹��S�h!�ʃƢ8)��0�#������6�W��.�O=��o���9��B�W�Ίx����(��S�4�L�X��0�\��hwS�܇������z�W��b4=I�����kY�u��X�㛃���rQ{�;�?�o���o�1G����T.����yp���v�k>m��=������i��l�>��k��"�9?��1>m$�\OK��Q{[�����qܪtƿ	�o�!�g��mޘ:j/�����p\p���Y������K��Y�:�Π>��e����]�+��eL�~�滎څ���G�s2���0�Ɨ�"Y���ߟ<o3}��ew�>ωn��D7�ӱݤr?���f�#�]��w?��L4���z����~���؞ ��_�	�S��|Y��g���~>|$ȿΞ�pMQ~����Vi�H�����kB���J;9.W�bϔ����gA�b���J�^�,����n�Ԃc�s=~OhK<	�g�i�/��y@g�_W��2�I��q��N0|=�[6����}��nً�S�q㽐��j>���u��������m�g]|�h��LQ�3����0뇗��G]뭶�#��z�t0�ј���Q�{�1^���c�_�Z��"+�T�,����tP�V������߷��j>� N	������d�����>�G3��Œϓ����S#�;�q��U�Jn�o���{.X^2�d�m7�S��g�1E����}ƛߞ�_�x�֝lq�sX�2}��=�/�q?#�3�/�L��"��mj�'q���C��S�5�2��@�0?���Շ����g�O��p������:�q]��v2��fq���}g���;d���5Ҧ������������_Lt��b�c�lS�:b|�ry��lt�-����ZL�cu����O�ϗQ~���^W�ԗ�������؎}j�:��Z�3A�qn}���ח작��<�~�{4oَ������HG{��v�,�c�ZD���+���n���Cl_�ܙ_�z����s��d���ιZ�l��m��c�����g�/d�Z�u����f�_������}���9§%�iշY}��Y\�����?���x_9�����o��Z�?���*���Ub;�(��h����������]����s�g�b���j�>�o[��n@���J�����'�CKY���d|O�~�z��C�#�ϑ_.�kw���2^w�����m3�`e�9��Y<W������IY����w�.w^�^'c;�~�c�6�Α^�֯V{���=�z�q�غ���\��a=#}��T�#�����Կ$I~��z���r�p�G����Y|l֫fg+��=#�����sf�d�d惴���?�U9Q=��4�/��ty��\���2���|�z�����r�8�Y���G�_�ev�u���:#+\����&៭�\�(���Tu��?.~>�G���?�y+ӟV���h�[>����WZG���|خ��٥�.���ӛ�D��-�sg����u���i�:��ds���C>S�t���ۚj��*�6+��ŇY���s���θ�3[�O�_�����x|Y}�J�~���"}u��8`lo�W��&��z�v�Ot���7���?�"N,�#-纀�����|��qb��]X�I(���ە��3-~]ܧ���6��6������9���u2�V��~�6��z�zþ�r���:�p_���'�D�ʻk�O$������\R�:��õ5�k�`~.�D}���S�c��ٰ����>�����ϣ�B�m�u��[Zw����L�?✑>�_5^F���|��a\�Y���8i��m#{��)����!?ƕ�����O��~P���z'�ŏw4�������[�y��JרA��R{N���q��)��[�y�ɑ�\�n!�1l�����T��Z$_�[�i6Ѷ���V�ͫjޯ��>|I�w��r����F]��"~�XZ�s+=��ٹ�Q�!����w���h��~X����3�F��pk����[qy��,�<��6��r����d�/�O2=O,��!�O"� �:5�}��z>��N��!����i���������ٽ0�c��ꏲy,����+Տ�Q>���(�W>?*��ƕ>+�휿��8O�P�3}Xt�y�R>��d�)��'/�}�z��A~�m��������ף݋������Q����ᓧ�E�{gQ��qD���a����q�o�_�������+nC��8�V��Z=.j����,�S~E�c���A>8O6k�:��B?<�]�u�7r��_��'���o,YU��Z��sI? �#���}�\����$���G�"�������P���p������ԃ���k{�:��_���x\��\D�����a�)�p�-�Ӟ#:~͇�?���9پ���sh��3����9��ܙ~�$�:Bd'd��	E/����g��u���Q$/��l��k��}���X��^Vw;0��U����.�'���QZ����H��t��k�O�JF�������ܭ���Y����%?���o��#���1%�]�m���?���$�V��9O��c�i���|-��[qqY=3�nY���Q�B�]����e���E�/���F����『v�Ѡ>V'�+>M�N}/� =�d��s^���t�G��I|/X�i����ܟ�\V�:�/i�^��HV�O�����B����v�bYU��S�t6(��Ǭ�v?"��36�G����+�wo��������,�R�k�qlgZ�5��%N�%n��+=�D�o�>��l�[����,5N����ď���ym�����7��WOV��d,���cf��R~����^�>语y;��7������L��W��[�#��/��6:�3��f�gM���45O,q�=��^,����{����ST������/:�����h��r�g�:_�C�̯��Wx^i�W�[@W;�b�⹿���]��)��#��Yʾ��y��`?��+-ҫB|�-=�,Y�91�K��Zb���J�pSٸp~�S�/�-�����Ι���fJ�����\�q�����r�~Ο�h�W�^LW.�g/+�_(+������=����+��y=5��⊴���=��[�4��eRO̯��X}��d�s$�ϭl��,N,�����i*߈����������p���;,���T�G�g�O~�4�w���y�<^h��0���M�h��^�CO@�x���g!�d__q\ěe��!��oyP���?v8�ߺ�~J�e�
�c�:-��S��̟�r:�c��ٓY�q��|Y��C��(����T?������ke�@|��A���6[����X���&חK�N��T��>-~-�!����h��wR����.���Rv�ᨌ��*�W���g8�9��?�ʸ�n�����s�#���o��G�vY=�DG}釙�������κ}��-��)y��ü�b������'������t����u����C�Y��vߏ�~ḸVW��e�iS.��:��Z=om��I�s*;�?H?YH��w�� ���3��f��/��ǖ��ڥ�᫹�6��^�g~��=i���ɕ�r�?������o�{��4�?D�h���<�s�������u2�kg���>�2�$�b����<��:���x�_�&�;�e{���� 뾩�v�~���G���n^����h�wH��d���]�ϞS~�s��Oĭe�������`�<G���镗�Ӕ>T_��嗖?|��ڜge�s�A��z���u_��2�@+NL�����B}AC��9�*�O�{ٸ�طH7;��#p� }&��B�څ�����ۅ���G����1�{����=�𚕽��/�����������c����r�\��q�~h8'�x˪��z�������{�����+d�6D8U���G�xB�������ֵ���q������Zi�kў����l�b����׵R�&�gP�z���.j�3�j]t\.��`�丣Z�5?@��nd��q�1E���BY�7TN�Z�~�N�G ��-_T�����
��5�I���v����p��c���Q��:�/�j>�g���?Ӳ������;ŏ��j��<�����{<71����t�z~-υ�>��u�Y|ޤ�v3?�Q��v�d�Y=�	��:8��������}�>��ov���qQ�<�g���ln�xE�I[�����ѿ�{7ѳ}nVOK��U�Ay\�]��;e5���_(V���������'�[����i�z �k����Ơ�,��X~m?��B|�����1�fx-n�ѯ!>sh�K���T�
�W=�:����iy\����|F�t^�/��>��/��/�2���j�#2�a"��t>�]��&�'s��sO��p����(�n!;�A�.��Gv����d5�>wܮ�?��nxIP.�D}�]��/#���#�s%^/�������:��΢΋%���uQ{�����)�S���fY��A��x��9�O����~���|�Y��?&~�x�h����L����7M$G�7��J{������s�Kd�0�F���6õf�]����w��6����g�^-L�z���3ņ>7��_��iy�{F�q�6N��S��VW�ٙ3��e��:��}��}dX��w�=[/���m��Y܃CT��+��1��o6���'�;ѹ��.�K������>fq�p�헏���qn��y��j~�ل�*!>����홻곾�����"{F˟��r�O����Q���g���[(���G��t�?�o�D����o��{ͣ�xb<1,w�t+;jo$GL�����q��?����O4�����D�c����8�ˈ��i>_��A[��g��W�?��5?�:�m���֣L?g�)�?S�P�_.�o���}Iӏ�9�&�3`���c?��w4?��ʲ��e�G�)�'ޟE��gG�uo���W�5�Ov��ۅ�@����zj�gT:�i���Q=��!m��1\�Y���G؟����^�;����r-���m}������l�3��D���C�:�`��K!�}���X�����.�������6d<^X�h?h���j=e{��ekM}">B|�4�C�@?�_⬬t����Ḹ�x=��g�J\�s�����X���y҆�0�����UV����A~��u��ޜ�o�s�(�����*V�˨\\ˣ��p@g<�&<ý�C7�0��t9�W�A�m仃~8��u�1��o�X�X\Xi��D�ds���u����E�=��b~{�.�'�ox����<7���|��wF��E{���b��H��7�!��C���岲?_
t��~�)}��ҹ}e-�kЎ��4��%	=�wܯE���ׄ�>�G��;H��{,��j,V+��<�`�=D��>�G;�
Iu�'�*E�mCb������=�sZ�H�B~��g�8Ƭ\�g��s��޿���y�$|��[�$����:�5�N�~x������ؾ~^+c�Ƒ���V��,�۾�����e��sԟ�+]e�?��x�]H����5�c�9$mqrl�g�eu��O�3�"�#�~;K�c�R�����U���L�^��~�����d�^Xb��h��:c���|E��z��S�WD���%�'���%��m,��q�H���{��#zd�d~���9:���g��ߟܮ��f�e~~�'�>�n�����c���a���j����[j��l���Bmv��x�v��d��p�gz賟�Ϻ�gI=Q.l}�r��g�:�'E�i��������n�fr�t�'�]�ԇ2��+T�ϣ:Cu�w&�A��L�=7�U�_��(]��_�N��N�G /��t�����v��E�p�?y��?�G��[I�qg���ۚ��`�T_�x������3&�{���e�W�?Q�+�����<9B�]}/:��ߙ�ߢ���ϓv�}��I����.Ï�J��{��7S���y�_w��b/a=��|/���{���=����u�눽�@��c��nA$>?��-��f���zm�E�'�~}~���j��K�e��5���'��/�w/��y1�iK�,q�ٹ���xu��iԟI?Ͼ��>���8Y��Q]�><O>���ϬS멥�D����6�I����!�������m����9��z����yP�m�:�U�A�׾�z�yMWg�Ͳ'�_S��E|���gp�n����F��M��s��ϟh?���g{���J���%˳���>;���_)���q��/Z��m��c������n�_w��|�포г�\O��*�MY�<��C�Y>�S���Go����h~�qDS�G$�����J�qC;$��7A�?-��pfW�+j]�^�f�;�����!�����!�[��������5�:Z�d6^���#<9���Wo����Y���|'[ǳ�ZStӉ��8�q���}S�O�?��Z��{O�-�8jO)��k5��NByQ�kw����/�_�;�C����A~>w�d}h�o(?�����˵sb�{�fF��?5�}�c�Z�vcd�p�T�隺)c=�����b�=���ײ_ԟ��͟s%>��5X��o2|��z�����w�?�E�3���
2�4淸E���:�OW:��D���ied��������.?��e�v�>��q�e��T}��S��,.�kqAu=�~��O���{�s������[b������G���O���7�g^w����U�Lu���Ϸ,>^v��C	�7y>Et���G$Ƴ}��&���x�h��}���U������g�
x���:�Q�d�߭�?����۪gN������ԟ\t��N�&K���ve8O����2�/��:�$�o׊w��S�Tf?[����x��~8S��=�{�z����i\�C	���5t�o�L�6�k��ݘ>���a��޻D�������c�ᬽ��>��qh�;�GJ���E����C;��#����T��|�e��%������e����xA;5��h�)V���.�-`��)Z�y��z�i�1]�������f��e��yn�g���sMmPݯ��ō��9[p�-z,�gq��~_����:��)mгu���y�FR�l]���CW�	t��h\�2Z�S����Ւ��Y�"�W<�?����xq����L�����l���d��ǽ�xo7�KH7}��3���J�:G�6*7�?p}-ϳ�7�w�!�3��ӯ��߾.NH��0�!��h����#�������{mo˼���>H���>c?�<�pz���:;$��:{/��V�'��)����PB�_���;
+�o�O�r����d���wo�tNc�r�o�l���^�M��6g��rq��uG{�J����?�������'������ɻ�Cn��J�g���w�h��ה�?-~|��5��ٗ�rF��O��0��]��Mn�?��l�}��}gQ�g=�����x|Ng�y��z)�c���������O�-�|���<�y��m*}9+{���@~��u|�W�7ֺ�l!����zd}���՘�5������T��*�%+<�˲�#Z_�����u�.*O'ď�xh�޳���i�����~��I�7��Y�A��g6^�W�O=u5��y��&�#��s�;�tM}�~`��W���~���b�|}�^>��xYS�g��ھ�ڤ>*g��XϜ����x��u\�j���� ?��8x>��k<�R|�����x�ke�#c2�a��ou��k�gq3,q<L�g�9�b7�躾�������h��x~N������oV�����]l�X�����+(���3�?�����L���sa��b��{���$�!�Q�.k��Q�TV�}Z����}�����j�W��L?��Tl�=��9�ۖ�?*�4�N���������ͤx���/�'>��,�.ۍx��E�����������v}��-���q��Y�=/m�;0������r�
��8m�e���a]��FF��ٍ��h�!�˘�#��3K�.�-�>������E���<�_F�CyGy)�ꞎ���	V6��l K��]���9|��o��)=��'�+�n�J<.�#��o�u��s���f�"۫����j�{���������hr��[p=m�;���X�Y?O'�#����u������56����R�~8h�7�?cu��o��_坕%��Aϻ[�c	� ���E�^K<ϱ>��a{;+��%���~�>�����G�e���������9P_�|S�Ӭ#�&Շ�>���+c?���?S�.H��ظ_-c}n�������//�~�4�w���!�E�w�����c��NQ},e��V��wZΛ�y.�c�/����'�o�����6���oZ֗d�=��\P�~!����>y�聬>�X�G$�ϲ?牕~V������,�_%{�zg���l]��ؠ^����R~��#ϵ�{+����s}�ŕE:�#��X��s|�Y��w,��b7H>��}��b�e��a�|U�oJ۹����S�;��x���S�{r7+������zN��3���V�ۻ'�w�seJ|g�,6��_�ٞ���{�z�G��@��5��l�"�:��"�s�od��J�CV�_��[f�V��ZiS��9	���8Ƭ�������\}j}��2�p��s<�Ð?���8���'�>v���ϧ,F�G�=���K�q�iY��U�����EվTߴ��W]�;����]�g�?�7f?Z����q�m��1��^R��G���gTz7U��D�_���5�=K���F�ٍ����S���'�[�{�}�/���)�?Y�/�E��~��-�C��R��%�{T��l�O�?�S����%[�3���%��s?�}�ߞT�9t;��u<ÓX�~��ӳ{W˝�)�����qY�&c{��A������{�>�7�gؿ��Z.ǽ����_Ge��(���Ey�z��o�χ���g���0ٷp�f���Keu6���}A~��\O�E�N@��e=�P��{�����8.8?��'��������[��G�=���	���U~� ?�Q�Q��y��^��o����D���5�?��t��I�?�gC�տ���SA~���k.��\��|�o[���@��']+m��)������u�Y�A-�����S��O$3J��>k#^��_�;�_ouB�����~�D��p����K��������'�I�'��|{C}��]�S���.������?Q\\��erqK}n�W�����5�k��\��FV�ޕ�����=%G�h�[hIe(�W.=��&�aȏ����s�����<b�Z��l��<���F���@㻇w}a��{WQ��l�nb��V�:�#��q��ɵ�8��o���5��pȗ�����T�гs(L��"�<�G|��[K�Y~�!������z�XE�g�o�2���/�۳'��/��n�����B:ڟxow^�!�S�V2?���42�� ��֤(�\b��~l�g�?YL�%�'W�������=�?@VO|���y�%��S�Z�S���*>���Ɖ� 6N:��/6>�(�%��cz���P��3ͧ6�74��������s�>#q)�o7J;}n)�<~m#���<����|�d�~$M�Ή$�/DG�s4������4��>k? >���ݯ�uJ��e�����/�e蝖��Օ�-��E�����*-��W�e���_�p �g��J��ڟٹ^v��������`�~�����'���Z��Q���v麠��e|����w����g��!��Y\�KeS�|z/`j�e>��b��e�e�r�V��ۼ!?�?�_��E���{��E���T���g�_y�7����������0\���h�c|]�W`�l-e��o��9����k�V܎&�u�C�1�٘s�u��iY��'�S�gʾ�t������Y}	h?�\�~�tP�����ø;�7)�\�@��s�V�_f�i��2?��5ܟ����~6oՏQ-�Ve��2�&��΃��������8�1��硶._&y\t����{%��:����2};'�ͫM��~��uޗ؎�������҆˲��cDg>���]�9�;!�1�=��FqV-�|8�Er=��s6i��4��Tߠ}��U�+�ߗ$	�]:�jw<L��Z'_-�*�wQ~��y���?���q�sL��}�h_pи���ګ�6��h\������Y��+[���d�r�x\��OTn��j��Y�_w|�]�����!�?��|��e~ψ����d�f�������J������]X��_@������+q<�;G�5�o��*�'�{����-�}sk�T?g�9;���D�3;9��.�ad��K��3���7�WJ�Ϸߠ�Q]��8��S�����������_���7=��¹��d�$�@?\��R�7�f�ma��1^l����G�?��q�Z����?����7$>�����]vN�r�O6%׷�:���]���/�t�_��>)7�cG�'H�j���u^#NF�p���y���}�%�W�C:���:��;�7o���C��6�����o��yэ���ѹm�X��k��<��Ծ��/�4��l������2��p�i�#�7��H7���8�(.Mf�fz��Y|�)���7J����7[��P�OK�<��a?��C��6��Q�}���N��_�=��,�����ʌ�����,�hd/m�z����Rݐ��[Ή,���5Ve4��,/vn��E��5��Ǔ���\K���SVwRY��T?�X?���Y��[���m��D����Xm|/$�٢xw�P{o����%����6���Ż���f+D�`dE����rg2��g0�E;y��W��{��S��-3��U�.J�./������▴Կ���qѽ��gt���o�A��������;�p>G瞙��y�n����7֫�n������a}�}�zY�=<Ŕ�kZ�gf�f�6#~S���uD������c������?������N[w�**7[���j�����]}@|��'�~����	x_�Y��I��K�^�33�W�ٽ�����+���J�OZ�%�c���������r��q��q�7OȾ/����)Ο�'S��s��	���O�����-YO���߇�"���������Tܿľ=�г����� q�p��_�W�̟�I=��=ڗev������{VV{�Hf�~O�A=��f������M�/�c�W��:�G��#^7Z�mݛ��2�S�fz��\�����]��#Ѻ�|W����u![w�����/��Ϗ"�v��x��]�A�cA�x�C=��s�m�{H�{UWHl�e�f���֟>�햩�{L���A?<��_��� t���vO\�|�A~�cf����o=Ǵ�j'`j�s2=���s�O������ݳ$���W�ߔ�w���+���x����Z�^V.��{dO��6��^W�����P��<_�W���e��ϗ��.S%�ǵ���tG{ǒ�u�Sx��շ�y^ �k��ߢve�+I�g����c\��>(���^d�o��e���d��t.��s�K蘟�/��]���Fv~�~3�x���g|�T�q=����r��8^�.�	�V=��F��Xd?���y��'��OߋA���I��}"�� ��틣u�uN�Ǹ\�+�t�Osi;��"�[j�7mv>����K���>��0�o����Ḑ~��z���:�V���A��o���R6">��<���gq\5�^���R�����B����̎5����<�����:Ǵ:��*M��-(w.����}@�l��~�ҵ����k~�R?<�ҟMt�wG�~P=���u��fH���H�i�]�23eWL�9�W?KV�q�^���*�ط�3e�}MPO�o�f�>���p�|N��8�/�E�=��oe�·V��ک�({��@79R�%N����O懌�?���^m��q��Q-�<�/���ϕ4���Z�5�a�B.7�������1��:\��Z�r� ��9����7�_t��8ƈ7��f�\ �zy��g���g��T����Ծ�ۋ�ك������Y����Ώsz֮�}%��y��OF�?���m��'$���	O��,^e��?G��-���)�<f����8�_�u�;�w1�����OP[	�\׃�[	����(��y@���q�������%w��O+���������~�xS�o�+�������oY}L�x�`��5l~������9�S�TwJ��._�3�st���X=Z��?'��[�y�x�g��ﻀ�ݧ��s{��Cٿ��-�cg��[����k�f�+�/H������9?��	��γ��ooY/2��8��:���*o�?o�ϝ3�c��X��h��k[��^�]i�Ib#ˋ������e�t�F�[m�W�^o�'���W����gvQ�o��e�������&���gvc�=JkWv/��g��ޛR>7~����U� z��/A~�Gq;3;9�������ge�u�U���7��O���x����i���!��_gG�ؙY���Y^ ��brv�&w�_��<��X���yS$/O��M��7�ON��u� �=��WZ~��5N�[d,�'j�{�c�����A�o�l/e�ݔ���r�����u���r�vٜ�v���B{��t{����qSYG�����U헻���jt{����U�o��z�|�8!*���MS~K��2�~���C�zϵa���������y��#F^��������of�L�������hm���8��g�ʵ��Sѹ� �ߋ�9�o����s��s��`�ʵ�v=�����~��g~�TڟJ�N�����}��u:)7��o�H<�y�����Sp�"�֧��d���f����o�������zϒ�9���x��]f���N�ȗ��w�5�ױZ���a��:nu��O��.o��e)�Ǳ>����L!�����a�S��c~;���e1��dr�~��>W6ϑO�c�>�|�������u��V6�[�L����^��ʝ��3�/��![��Q}2<@�z����:�O�Q�45��^�K��۲;���t��}�F�?;��}7��cm�]f2N	�w��������7�3�ʺzb?�~��8��;A����:�-�dĉm��$�R~,�"�/s�q�:�����$�3|Z�w��/Z�l���߳t���x�P|\�������I����Z�qp=��Y�gj����=�O���f~`K�����+����9 �ʘ*�ҹǻ��Dq=#�Wu�_c�2����߲��G|�ů��md�Yb�7��g~	mǮ���0�~0�+��������w$�Z>}�&]? q��,n�>_���=\��}��������7�����d�D��<?�8��Z�Q��4�g��3���w;���S���q����H���eD�sYi��}%�oy��mh�KZ�ȯ�nݏ�e��� ���a����+���^���mgt����9��de`��o�~���'�D���1�Sdi�������(�>��d޿�x�;/n���:V8?�}:�� v8�{q�_�5V�����_8Lt��E�2�_g׽�~����a܆)x6^��������Qj����y�����&���S��,~��}+Y{�����>J�֩��h�ω��zM�b����Rf��Џ���~�v�]�|��u.#�
ۊ|p�����8�!���℞�G�?��(�:>����E[�����������9�%�D����?(����O�|���Hޣr�w������L�V���z���jK���?�4�{�+�
xn)�̷\��⌙��x	���xVF'mr�m���������>Z��\��{Q��{X�7��`{�]�g�~-�m�8���u��{��E�v����$Y�Y�cL�~�za|���������Q��Y��u����t���/��)}��V�� ��A�g�㦶�C�슬]$�d�\qG�Z������<��S�(������pݹI�?p�>N��G��������gtK���u�J8�Q�0f?���.8��Ƕ�3{���--vH�Ho�;�m9�g��~��Γ��w�L������ǯ��*�����pd���Gv�LҮ��?UF#lk\wK�6|�%	}J��u0�?�����#�g"�������=�7���3�R�o�4E_�O��y������8tm�S��'��=�e�U��2�&��d�>����/��WO
�k��!��<io��d?�c*�����~Q����)2�y�����h?�|�O�gwx�	�aJ.Z�#�N?�����ҧ�S�rE�������o��s4(�]��_q�<%k��.���33���l>O������L�Ǔrq^�;߼D��;�_��=�����I.GX�Ϫ��e���"��Fg\qVnv�!I~l�2�����8y�U�3��<�ۼg��V��� 3����Q?�>�nj>����Z5��t����9�jf�9��O���<| ѭW��S���3�o6�to�����k.YÇ��|S�?@�<������~^�jߡ��[��6���>��l��ٙYgg��x�:8{n}>%�{�v���R�Ą�2���������N6��A�5��Ú^{�g�m'd�>��z�9E˺`���,�7G��W����a]2?��[������7����3O��!>S�"�STn�����W#���t���?�oM~bE�M��x�C!�^�/�v�? ��e�|�|��B|c�Q{�ss{���|�����W��M�O���*��r0����Ю�Ν3��k��4<��k���V�js��T��	���#���ݢu���㠭���Y�J?��:��J�?��j�^^>��a��$A�V�By��)���!��h�e�E�j�7������r/��|��sk�Y���Ƌ�S���:]��x������y�����-;W����Y�n�U.��yb_q�������x�BY=-�½DW|í���%���op߁�)lo�T�������?��-[���y񞑎�+j���L.���"�~�0�[��)��i��U����S��ٙ��[�H�y��W��lO���a=lkg�g{p�������uvcfo`}���x���q��=��[�@���/��b>�_����JS���M���n&:⽣}�����(��s�c�ly�S���2�35��>g�￑�L�W�u�\��?¥����v�ɚ�
�o{S��UO�>�*��A��z�z\ϩ�?��U��S��oo�C�~��X��f���ӕ6H����a��{a\.���?���ou:Y�棸f|�����ݬ�}�\���j��sd�s��/���Z��)���?�G����"~]���G�=feD�2�ɦ���^��D�m�:e�F$�x1��şM�+[���#���?�w���g��?!������W�|��1�0����f_^G���q�,ݟ��|2��R���]������JS?��~My�[�g�$������+�� �W�6���>�r�|NǍ�^Y��K��J���f��q��d_7F����-���{.��?N�m�3n�F��<(�Ub|f���m���QH������������'{��%��S���u}��gqH��W�l��e��ɵ�2-�w���{��_T��#��G���7���3}����F$�7-� ����H�)��7�է5����gx�u��nzR����z�o:H�=�����c��[�/��u-�T���|�{���f���M�Ο�8`�]d錌����[a��Q���O����nG><���Y<�V�Ɣ�~3E�*7��������-�m���#]�Z�]"�8`�Z���ˌ���d�)ѹ��R��2����.�/�]�����se<ߦ��lg��O����=,��<A�h�>�'�#��~�ijl��̎�x4&�������C4Z�I��!�?�A���e�y}Z�?N����y#=�æ7t���w;��fh=��D��<m��b�_"�X�F���H@��W�ꇷds����Լڦ��5!�7;�@���޿ 	������Q�(�L���wʵ���}�5���G�5�N��s��8Ȼ��W��ƺ��f���;��X�����*�t�D�	�o���wb`�X���$޿|H��-���~�ˈ�ů��g�(�>��X_�{�q������ɥK�Q�����o/S���F�'�?+hW���R&�,/���2=�>O�pD��S4���|�cz���\*�y��CV�'��U�跖�/�=������Sd낽ϓ�no_��<έ��g���O䝝�d�n�ٓ��,G*�W�2/����\l��xa=��n����>:��Z���5��8��sZ���qQL�����x�~6��?UO<����m������Y���y��?���jWp}4��G������-Yͩ'�9~)���j�F�i6�������%���bv�����L����p5��3�?!�W�����5��E�!>>���O>"{���г�����'�y�?{/��L����l?�}��'���g�gX���b�\V�2����Gd�ox>�k�9#����}7��,?���A�M�� �ؖ�ވY�����~�v�]������:����~��������5�e|-��A;?���<f�[����|�?�Q�.�{|y�����c��?G=����VQ�6>�79��j�\d��o|��?9��'[�'d��z@y|���n��7���̎j���ڍf�_�N"�geD����8o��vY���%|Zޟ���ZZw�����\�Bɦ������k�n�a��Ծ8/�cg@���i�ox�"��>A��'��Q�x�0=���Uv~[V�_�a�������x��l�7�=��t�8����~��9�'���|v���ϟ/�-�+��=����Zby1��A���oSm����3<W&w���Ε��G��W���0������'�l���^W�A�oV{�pԭzuʟ���~��~OC=�~���1}�|0�#1.�~��?t�u�#�9;ʑ�}�C���޻��#�q? �\My9�ek�/A��ol�r�b=�2�c@߬4��A�W<�w��$�{�G�xQ|?M�)�'G�.���`j�G�v��e�x�:��]v�h�6�[Y��w]?���Zq��>\��@�q��"���y������u���oغ~���e���ƽa�R�jK��Lٿd���"z����z��#|�:�1�;d���u������^b��bzv��������誻n��~0��{�5���~C����\b�����3�Ù���G�x�0Zn<�o�yٯ�nY�纥��%������nn�i}M���{P�։J3�K�^��Ώ�R����"����z��ŹR�?[�v����ה����o�u���t8�t=��	�	-e�g��*Dvf�}��㷣���o����9(��u�����L?p?[}n*ED��چ�{����ݑW�s��߰W����P���񌻟�ćo������q�>�W{���蹣灞����z��;���n���G�zjOO��{z���T~O��Ԟ��T߁~?��T��wA�T�����ئ��&~���m�M��&�K���꿤�T���_R�Kjߒ곤�ܡ��P}v�>;T�����C��p��?�T�]*��۵ߟo�y�	[L虰`�6���3�O��#��c�O��#pM;.���'��\=��z�X���=ף�bn��<�1p��)�e�U_p�n˂��z,�����6�d��a����U��R�\�%�t��.��%wᒋ����Rv��.e���ʎ��c���vL�00a��%v��c��X��-��W�e���fW��A�ʠceб2�Xt,��~ǲ߱ w=�i�m�)�z7p�Y���K�b,�Kvǒݱdw.e�mYp[X��m.�e�c�ﶹ��%�cA�X�;�n�5��RX�;�n�'���å���r��<.�.�]j\�ʠgeг��,�=�~ϲ߳��,�=Kv�ť�d�,�=Kvϒݳ �����ܳ ����=˫zϫz�ʠgeг2�y��{�k���C�ڡgC�geг2�Y����,�=�zϢ���osMY��zV=[=[��[���g�ѳeгB�Y��K�k��5L϶C�*�gۡ��bY���rzV9=k�~�����:��Ų�2��2�RX)l����Rk�����Zj`e`�5��1��c�b����R����폁���zl`e`�6��X)��VJ[(���e4��BX)�؆� X)�V9+�����c����
eXr)�.���e�aln,�����?��lL,�����?��d�r�`�]��.�#�`1]��.ؘX�1�`!\�.X�,/6l,x�_�`[�`�Z�2�`[��~���Ђh����h�&����/�^�,s^���/X*,�^�,���K傗���W��������o,������&,X�,��m^��yE�fA�fA�fA�f��f1���t��v�7ۼ�n�do���k�6��6��6K�6���,��,��l�o�J��+�6/|�,��,��,��,��l�o� o� o�Z���LYn�YL�YL�y��f1�f1�fk|���m�m6��y5�fKz���m��m�m^	�y��V�96��l�.Y�,bK^+�l�.Y��c[�T.Y*�,�K6z���.٤]�T.٤]��.YL�l�.Yn��D/Y��,�K^���f/�
^��/yE^��/y�^�ѻd�_��/Yԗ,�K�%��K^՗,�K^ė,�K^o�,�K^M�,�K�%���tɋ��v�k���%K��y�&�y�r�Ë���/�;,�;,�;,�;l�d� ��j�Â�����������K��+wX�v�,�a��a����v�en�en�en������^owX�vxy�a�y���^owx��a1��x��v��^�w�p�aQ��%z�-�V;�vX�2�a[{�m�V;lkﰭ���c���;lZ���aC`��+�V(��PvY��B�e��˦�.k�]����e��f�m�]V9�l;��e��.+�]�.vY)�R�e�b���.����v�2�e���:h�u�.����f���+�.+�]�E�2�eQ�e��e��eA�eA���.�.��.��.��.��.K�./⻼��T��{��]�"l��oǻO�e�(ێ�t�Gq�o���\Y[�ϖ�ӹVt��}²Oqeu�]�kW��s���Oq����ޕջ�z����5���gu�S\�+k��,\�-��p��p��v�/]�K�y�zl����v\��v�x�V�8λ����8�V�V�ҝ�n99݇��Sx����n9��r���=ۧ��lm9>Nr���n9��r���$w��Oq�q���dy���>v�>��������>~m���r���dykp��,���)�N��qk���N޷�W�W��om��n��l��l��l��l���v��t�;M��4ɖ�$[N�l9M��4�>�m���r�e��-�[�v]����u�;����ϖ�6��}
קs�s��s�D��O��O�,�}��>�q��vNGuNG���)��N#uN#uN#uN�tN�tN�t�+���Y��%:�:�[�at��+7�.�m:�m:�m:�m:g]tN�t���&�&�&���S\:M�-g�tN��c��)�W���n���S\}���m�9+�s��sZ�sVJ��F��F��F��F�,���-������+��8z�Iz�Iz�7z�z�zgo�N�N�Nr{�蝝�;��w~�d�w��;����NN{'��[�{'�����Ie�����i���v�r��/]}��>N�{'˽���Y����In�$wڶOq-u��;ˡw��;��t�N�{'݃���I��{pV��{��Oq|��NN�vNr'��[�����ap�=8��J=�uyp�>����4��V��������)�>NKn������j>��|p������/���������n�n��bp�fp�fp�ep�ep������)��?��%��gN�n�18M2�=��v��-��-�7No,�U�pzcᬂ��
n7�pv��i���,��Y8��p����o,��Y8��p���y*N�,�nb�v��X8�p6��i���Z��N#-�FZ8m�p�e�t���&N�,��X8-�p:a�,����%NK,��X8-�p6��i����%N,�X8�d�t��鄅�7�w�p��i���@No,��b���Nol;-��t¶��m��vҽ��	�N޷��`�����@���v`�i�mg]l;y�v��dy���7���n�Ƕ�%��d�Y�N���to;;a�� �N���,o;Y�v���$w�I�m��o;9�vr���t����Ϳ��k�K�[s�ݚ�����������[��N���_:��ҭ�K�R/�J�t+��I�ҭ�K'�K'�K�R/��a�vK'�K�/X�uy��t��t���[a�NN�n�]:�]:�]:�]�]��I��I��I�ҭ�Kg�/���t+��I����K'�K�OX��z��}���;�\:�t�t�t���Y�K��[��z�|K�v/�J�t+����K�./ݺ�t�f�4Ɏ�$;N��8-��Ď�;n5�qZb�i��O�qzc���v����Ď[�w���q�����8y�q�����8y�q�����'�;N�w���Ux�I��
�Ux�I厓����8ky������g�8��q�򎓸�.�8��q���k��׎[�w�j��dp��ஓ�]����|��鮓�]'��N�vݺ��l�]�R�:��uR��p�NNw����l�]���:��u���[�w�e����]���:�|�i�]�v��u`׭��n��uZb���w���u6������u{�]g��:�`�i�]�mv����Ϯ�6��*�u�f�� �N��:��묂]g���i�]�v���4Үۿ�:�`�Y�n����خ���:Ͷ�4ۮ�c�N�9�b�0���;��Q�����Q�C$��(�3k��a����:�Z�F�P\鬑:�H�"�P\YlotX(��k�Bq�`�S(�t�?��Jg�ԝe��9c�p��C-��[;�C6vgyWR(�7X#�S��
�ՇuT���`U(�>��:��,�R�H��L��3��a&;��,�c�[:���f�s��n�-�n�����f�Pg�7f�s��!$;��출�p���a&;�����s��Ρ�-�[:�l,�?N�8�c���؛�9<d���Ɩ�[N'8c���q��;�c���s8�Ρŕ���n����-�@�-�@�-'���m�-�9�b����vm�9�a�І��v��A��J�s(��s��v��S�,��I��v����I\�$Ρ;���ޯ�:�_�9i�x�P(��[s��sX��a�:�����sX��s2�9tx����:��+W�[Oޯ�TvN*;'��9�_�{�C�u�t��un���:�_��~]�d�s����C v����Vw辮w��;YvȽB�V8,_�;�v�Bq��5�wk��v�[�{�0t��n� ,��ޭ����;�`�;����CvI��npH�Bq�qv�Cv��m�9la�p�]�t�CvI�9�`�;yw�����ޭ�I�9$a琄�C	v%�����J�s(��! ;���ޯ�px�np����w�	�&�P\YN'8�`78yw��Ρ;��J���p���Jw6��v%�9�`�P���v�N'N8�`�0����! ;�����s�Ρ�:��+W��w���r�P\Yn�w��!�:���r�sȽnp:�a�������i���	���s�npZ�! ��rx��a�:���*�[8yw8����
ŕ�v��r�P\�NK8,_1�g�t�W(���NX8�0x���r+���u��9^�w��z�I���u;�9�\�8>N*N*��sh�n��t����������I��I�C�u_�94]��t��I�����s��Bqmw��0x���
�g��;��+n���l��~�|������V|��+�.'��n�w8�Bqe9��v��9�^��l�m'��N޷��|�C�u�n��vZ�a�:��+W��ޯ�v��m�[�P\�N�8t_�pzݶ�	�N'8,_��t�C��k��	�ί�0������w�,�cN�8la�p���v7�9�`�p���v�9`����Np(�Ρ;��&�P\}��X:;a�����	Kg'8$a琄��i�-�n�t�e�t�CvmX(�,�[��s�������?��-��q���!;�H,W�["�s�����qv������H��9Db�����v�-�n¡ŵ�韥�$[X(���I��sH�n�i��I��s������S�q:�a;� ,n�C ������}�I���)�8yw��n�i �6�ڰsh�Bq�;yw�����'���9Db��v9;a���
v��:�b�P��C-v;N���s��Ρ�'���9c��>t�����c,�
g]�8�¡��ֱs��Ρ;�Z�F��u��0�ݮ�F��u�î���s8���;�Z�v���uv��v[��:��І��j�t�������9�a����C�+�i �6�ڰsh�n����v�jݮ� I��:y�u����T8$a�8>N�w�J�P��C	v%��:�u��! ;� ��s�Bq=�g��Y� �C �X(��,e�Q����ò�;`��~�����׻x��C���W(�,�����.&a����wq{��n�wQ
{��w(�ޡ{� ��w��! ŵ�}�C �ػH��Y�$�����W(�]l����;,_����r���w{�����w{���N�P\}X���;,_�{�C��."b����׻�����;�_�ŶD�ŶD�0�����P�����;�`�P����.�a��������;�^�{�C���׻H���	��m�;�_��~���;`����[X(��k)�	��R�;�_��[�S��wq{�	��w��! {��w�{��w����?�]��~�m���?,�v�_�X(�,�m���r��E2�"�w����6,.�!����Q�;�7j�w��ޡ{�w�{�l���w�{۰P\��Jq���!{�l�]$þs���-���w�{��w����-�ֱwX��a{�u,�.�ֱw���E2�;�m��w�{����w��ޡ{�~�]����!{�w��!${���B�wɾ��M��v�;dc�b�.�aﰎ��[ػ(���R�;c�p�z>��j�w�þwr��.Ja߻݄�1���e�l�]l�����Y��;Db����;�a�;9u�þwR�"�mػH��C�m�;$a�P��C	�%ػ肅�9���U�E,��Ɏ��;�`�������w��! ��quv�58�r�{��J�w(��a{� �'_���'_%�;�`�P��C �.N`�0��C �.*`�0����.*`��7�;�`�P��C	�%ػ��C	�%�;`����;L`���C���W(�n�sx����z���]|�ޡ�����.�_�p�! {�w����	7ػ����W(�t�I��w��ޡ{�	��_8�p����]|���{��]|��!	{ͯwH��!	{��_8�p����.v_�Ⰵ��i �w��~�t����w1 {�Z���w��z�6���w���!	��� IػH}���I�;$a����;laﰅ���[�;laﰅ����NKl;-�������;�a�������N��肽�.�;�b�0���(�.�`�P���.�;c�p���.ػ肽�1�+�i�Z�"�w���!{�H�]���!{�H�"��v�a{�H췝�q�{�?��.���]�����"�l8�I"�w���!{�?���w��~��m�[��nq�{۰w��a{�Q�]���E)�]���a{�Q�"�w����$���w1	{�6���wQ
{�-���ph�ޡ{�6,�cnW�І���K�ڰwH���{��]$������ %X(��N�J�w(��E),�����%ػ(������n�w����-,Wg�8�a�І�C�.�a�"�Kg�8Db���C$��ػ�����/�FZ:�䐍�C6�.na����ػ����(�.na�0���(���;�b�0��C$���;laﰅ�C�;�ᰅ�C�IX(�t'�I�;$a���a{�-���wH����'�."b��,����w����{�?�w�Np���!��\���E_�j�w��~��$��;Db��1���;�b�b-���;�b�P�����;c�"+
�k�Y ��;�cﰎ��:���;�cﰎ����;�c����~�]���Eh�]���a&{����wx���!{���w�ݲ��"�wx�ޡ{}�wx��aŕ�4��C����:=��C?�.�b���C��ػ8�����;�d�����ػȊ��L�3Y(�]N��8���U�W�;\e���{#�ఎ�C6�88d�p����"".�����C."������8����{���p���U��΃CZi98����C9���C?�̓C?.F��b$�88�����8�����C9����CH.F��b$39�����8������88\��p��CQ.���������6��P����88\���+=���CZi98\��b$W98\��p��CQE98������CY(�.��Brp���WzpQqpo\��Bq|��p1���rp���a&��frp������\����(���rpq5qp����*G�P\YN�8��CQE98e�����18���𐃋�88�����C9���CH.����<��?398�������88���Џ�C?�8��?98<����C��υ�j�4�CH!9�����L39�7D�у�UWY(�,�m�����rp1$ŵ�����rp(���(��frp���a�qp�����Z�{���qօ{���Џ�C?���Irp#1rp���Ő\���(���rp(���!zpQ%�KwQ%���;�yrp���Ţbsp���E��sp��E�ܛ���ܻ�ŗ�Z�l���sp8��ū�sp,��\���!?�rpX��Ţ�{��^tp�*� �tp�)� ^tpx����zp,�)�tpo�ܛ��rpH��Ŵ\L���U�VZup���aS�rpQ.�_\���Ž,�N�9���ޗ=�h��C�.Z��e;8���g.~f���8=氲���+;8���"j.���г�C�=;8���г�C��M܅�z��QO;��ua;8�������98���0����.��P��C���܃���;8\��p�����;�x��C��;��u�;���{[�఻���9���{[�����.z��w�;84����=��u�k�Ӈ.�����C��;�7z�;����C��;84��м�{��м�C�.R�����..h����~�Exp��a��\���a����;tp��a���-��i���Z��\���a��r�P\�sX��a��
ܛ��F��� xp����xp��xpo�xp��a�_tp���!~���P\}��p����{��vwp����p��
wp��\4��!u��RwpH��!u��-W�� �;8\��p�����8:�w��;����A:�7�<�7�<���C�.��఻���.�����+���\�����
.�����-��Jq����2\,��!��tp8����tp���!~���wp�C��RwpH���Rwp�C��-n��&:8|���.������&:�h��� �;8����{�ࢉ�;8��ࢉ�;�ء��:�H��C�.R��0���:8�����C��m惋Z(�t�[����\�����tp����y���wph���y���wp�./�Rg�8|���C��;8���p������僋A:���{���"��;8�o�����q�K�Nxp8�Bq5t��C�+��-9<8��࢒���+�Y9\(�>No8���p�	.i��V8M��4�C]<�w�o<8t��ă�J:8t���ŃCK<8���pC<8T��P��� �;����C���1�������wp���!~��\���!~���wph��aw��vwp����K}ph��!u�v��aw�����:������C�.N�����{���ފ>�8��C�.*��p�����������?[w�#��k���3K�(���إ�1�>�Z���`ʱ��@?d�4�A�4��=��{��{м�;���tӃ�=d��x~p��{p��,�û�ɥ�w�'Y�I�i�{ߛ�ީp�ߞ���|*A�s���D�&�7Ѽ��M\n�r��$�&	���M�N���D�&�7I7M|o�{�t�D�&�7���M2Q�L�D'*8�DMTp�����$5���M�o�{���D�&)���
��ݥ$)��Npb�<��G%oEO�U��D�&�7�VMpb���{v�U���$[5q�I�j�����'*81�ɛ����$[5q¹�H8�$5qNY'���N��ӑ�ĉN�V�µ�[��(y{��K�X��'��.N,q�њ��$�5��IFk�o�$�&���7N2Z���$�5��������&J9���*QʉR�
��ᖓd�D2'�9�̉dN�_����6'o�O�`���Y>ȉ7N2Z���D 'o�OLrb���
�}���d����;��<��}9ɃM�t�(�D)'&91��[�sӣx�}�㚸�$�5q�IFk�ȚH�p]��s������-'n9qˉ[N�r�����$6��Sa=tlsb�ۜd�&�9qˉ[N�r����{���-'n9I�M�r▧¹�H���$O�s���$'9I��
+����]�X��'r8ɞM��T8��|��'�8�ĉ%Π���q℧ٷ��'�8��	'N8���M�o�s��� 'Y��
NTp�����D'81�S��Rpb���$A7Q�S������&�7��M|o�{��;�n"u������&.7q���M\n�rs���D�N���%��M�m"l����&�6��M�m�������&y�I^n�i+���D�&9�S��v�o���$�6����M�lbe��z�I���&�6�.A�n�g�¹xNA�&V6�����
k�l�`���D�&�u
��@nb\�T۩p>˨ש�f�/p���M�o;��3H�O��&26q���Ml�^����$�6q��zM�k�^��کp.: ���Mlb\�ש��U��T�.>�8���&6Q��zMk����ĸ&�5�I�m�a�d�&��zM�k�^��ĸN�뢓 Zњ$�&ɷ�qM�j�U��d�&�u*�Cv�}Y���Ml�|;�*݆�۩�^)z6I�M<m�g+�X�D�&�5ɰM�kb\�:�̮ �d�N���7P��zMrn�8�$�6����Ml�s���&�5Q��zM�k�^���$�v*��ɷI�m�`�,ܩpv�/����Mdl"c���D�&ɷ���
+�#���x���&y���M�rs���D�N��*��26��S�]!26�����M%�G=
���D�&26�ԝ
�k���xکp.:	��S�gAoA�&26�����
+�Ʌ�ݩp��5��M�k�����D�&�5Q��zM�o����d�&Y�S�n�%г�H�
� $�&	���M<m�iO�x�$A7񴉧Mt����&�6��M�mbna;��	��(�$A7q�S�\�n�p����J�n�ps���&
w�9�O�$�&�6���M�m"lO�xک�B��𴉞M�p��q�6d�&�6I�M�oO�x���&9�S��7��Mnbn/�v*A�P�T��������^\���^2u/
��p/	��{Q��{Q��{Q���o��(܋½��^\���^\�TX���E�^��E�^����^Rv/���i/����{Iٽd�^<���^�p�������^�q/��b\/���s{ɹ��׋q�׋q��֋h�hՋM���K��T~h�K��ů^��%��"Z/~��U/Z��U��u��ů^��E�^$�E�^��%���L/���a{q�wzI���Ӌ;�(Ӌ �ҋ �$�^�%���E/^��E/^��E/���</���</���</���</��:/��:��{.T��|�ɧ�΋ؼ�͋Ƽh̋Ƽh̋����^�_�������ˋ��Hˋ���ʋ��ɻ�|!$/ɮS��w�Sa�|*q�WyɃ�
��s���Hˋ��H�K��%W��+{��{y��iy��iy��S����iy��Wyq�3yI�ɋ��xȋ���Gf����LN���7P�EyɃ�(�K���U^\��UN�s���׋����^4�%��3/y��<ة�:y��9�L�Bc^4�%����zј�yј�yј���K��El^��%��b8/���zId�h̋Ɯ
k�o�\�Ƽ�ˋ���˩���yј�y�|�TX!O΋�΋ϼ�̋ϼ��Kj�ElNų���=�d׋�
g�G!?/���z���׋�
WAo�y^�%I�b8/)��9V���y1��y�D��͋ؼ��K&�%�b8/	��y��ԩp�ؓ�wz�;��ϋ����Q��yQ��yQ��y1��y��yI@�$�^P/��b8/���yQ�S��|�Q��y�=I��	��yI7��~�yq��yI.�
�bO��,�%�t*�����R�S��t��T���'��^��E�N��U�I�/zIR�
�Eo��^,�%�bA��{.�/zѡz���$�K��E�^2Q/�s*�.A&�E��KO@�^,�E~^��E~^��E~^�M/��ez�2��ϋ�
G�K\����N*��p^�%���A:Vȷ��΋꼨΋꼨΋�$�N��H7��ϋ���ϋ���ϋ����ّ��9��s�<����@~�G� I��C/��zII���A&�ł^,�E~^P痗s�I�/z��ԋ�xы�xѩ�B���/z�M��^L�%I��E/^��C�%p<��C/:���z�zѡS��=	٪/z�V�ҋ�XЋ�XЋ�΋�΋�Ωp�<��z���l�K��%[���:��bJ/����zQ�Az��ԋ�xы��Ћ�XЩp�M�L��
��nC��%u*\)�Y/���N/���zIm��өpv�HHԋD�$�^l�T8;}�zId��ԩ��6(�K��E�^��E�^��Ŕ^L�Ŕ^2Z�ңP�S�n�0�S�=���L/9�Sz1�SzIm��KF�ŋ^��ŋ^t�E�^R[/��S��Ϙҋ �ҩ��Y���׋2�d�N��LGj��A�^�`/y��<؋V��ԋM�Hԋ)��ҋ)��ҩpdvDM�A�^$�E�^�^��z�H��K��%����z�ezQ�S��q}(�G��Ý>��C�>�Ë>r\��:�ա�����|h�Gn�<������#I����HR}8χ�|8χ�|8χ�|8χ�|8χ�|$�>�T�����S����G��#[�����V}xч}$�N�;��Y~�҇)}�>�#7�aJ�¹~�n���L�t*�wl��.I���HR}HԇD�
��}�y�ԇM}�Է�?�ԩp����C�N��ӑ�S���(rS�¿���U��S�*�6�w��0���0���������HR}ש���u*܍�=�#I��`I�;���.�gz��gz��gi�SaͿO[��թ�f�!.��r
��p
w*����}(܇�}d�>\�#[������S��t�M�ܿOR�D֩pzv�awI���м��м�lթpv��w*��^�~�߷�u�G��T��:�W��S�gA�#��a���ᄧµ��7��
~���}�߇�}�>��#I�awv�aw����м���M}�އ���z�}�]�0���ԇ
~���|���>\��
��p��{�q�/�� l����������G��T82�\��C�>��C�>��#��!l��!l��!l��z� �.%ؓ�p��an����o���HR}$�>4��ow������lՇ�}h�G��C�>\���N��\H݇�}�ܩpv����iV��w�p�S��χ���}8؇��
��oW�;8؇��
k�K�e����,Ӈ�}d�>d�C�>d�;t d�#���n��\d�C�N��p]|�I7}�؇�}��>�ø>��ï>��Ý>��T~׌D}d�>l�C�>��TX���Sa=|�� ~��UZ��U�����NN�ï>��K��֩pv>ݤ�>�L���^~��U����S����W	����S�\�}G�>P�������H7}��>�M��!Z��!Z���Wy�����:��w���D��#��a\~��WZ��e��S���h�
g�/>��!Z���H7}�ש�:	y�;�Co!���e��2}��Gr�C�>��æ>l�æ>2H6�aSu*�Uv��ԇM�
g�`S��rJ��{d��C�N���)}�G�#q�aJ��!H��!H��!H��!H^��E:��&��/����|ѩp.>�x�G��Ë��� �Ї}XЇ}XЇ}X�Gv�Â>,�#;����������H�|�χ�|�χ�|�χ�|�χ�|8χ���
q�S���
p��4�G��TXO��>t�+�eH}x�G��ËN��g� }d�>��#)�aA�aA��$8�Gv�#)t*��P|���
?/��&�H}��G��T��b�@��C~>��#q�aA��A�С�С��ч}�χ�|8ϩp7�H$�>,�#q�aA��!?�����Gv�#;��:-������H�|�̇�|$|>��T~�3��(f�a&��S���9�(	�W�H�|$|>>��!-�r�xr.����*����p�W�p�W�P����G��T���Y�^��p�Ezg�*���"��H�JR�ȿO��,R7{Y��"�������M�?*����\dl���,Tg�:�9��O(�g�<{Y���^����,\e�(��?�
G��t��x}��Y�����,�e�������
����](�BQ��P��~,�,_��B?�/�c��XX�B6o�/Db!�Xdl�E�f��Y��"us*�?A�c���������c,c����B6��xG|��X���0��Q,�b��Y��BڰІ�6,$a�X���P��,�;7X���J�P��,�`���{v�`��B	J�P�S�\��>a�I���.�a�������?,�a�����m/Db!X�������Sa=�0��Q,�ba�X�B$"����?,�a�nZ��"��E�i�nZ��B-jq*���Z,�b�JZ����c,�K���"��H.-�c��X���1��p�����X����u,�_��B?�q*��>�u,RI�T��m�u,RI�T��C�𐅇,rJ���"���)-\e�*WY��"��H.-�KiYx���,2H!Y��C��E�h����B?��xk|a�X�Ʃpv�wH-Db�&Z�������?,rA����N�ŕ��%��0��Q,�ba�X�wjq*�1>��ɽ��,�c��Y��B6��H�,dc!�s�:)��~,�c!�X$|N�5�D-j�P�E�g��w���p�E�g��Y��J>�$|��x�{�n����E.ha&���"�xo{�*EY���Ly�Ezg�(!Y���~���2����,�c��Yx��C�p��Z,�b��Y$s�����=���x{!�X��B$"���,��TX�y'{a�X��B$�����$,ޜ^�eڰІ�-,�2mX�K�ІE�f��Y�K���,Db!�X��������?,26X��������6,�a�mX���H�,��^��(N�#�WG-Y���Ջ��"c�p�E~f��X�gj�P��Q,�2�X�����E~f���"Q�H�,dc!�X�]����u������:��ŻԋD��:��xsz�{Y8��1���l,d�T�.�ֱH�,c��X�\oE�
WA�:N���'�!�7��𐅇,<d��X�����u,�o^�����~,�ca�X�UF�0�E:e�EY��B-j�P��H,Db�`9�C��()��Z�
g�o��B-N�#�[p�E�e��X$X	�E�e!���"��ȫ,ޥ^$X�ȴ,�d�rY�\��H�,\e�rY��C�p��Z,�b!X�S"�����Xh�BڰȢ,�a�mX$Oɓ�?,�'�XdQY���̋t�"��xwya�t��:ֱȢ,�c!����m�Ee�!�X$OɓE�da&��ɩp���d�EY���LB�ЏE��T82;�c���U�� ��0���,�d��BQ��P���,�)W9VH��^oW/�e!-�L��^6Ҳ����l�*Wٸ��U6o<o�x��^6�ј��l4f�1���7i���l�f�3����Fc6������l\e��٤e6٘M6�T8�o�i�f#6�����g6o<o�f��و�Fl6>s*��4>���l�f�3�l�Fl6b����֛l�Fu6	���l�*�7�7oNo|f�3�٤S6b�I�lޜި����M:e�EټK�q���l�g�<���w ��l�g#?��8�&�I�l,�T8=����F~6γI���)���;γq���l�g�<�t�&�����m,h�3��L6:�ѡM�d�E/�x�^t�!���O��8X�Ƃ6���M>d#?���Ƃ6���Mbd�<��8���M�d#?�µӣ��M�d#?�����y6�s*\��w)��l�����g6>�ј͛�Wٸ��U6f�1���l�߼#�y#|����&��q���l\e�*Wٸ�FQ6��Q���l2$��&1�Q���l�d����pdzB��~l�߼�ɇl���x�&����l<d�!��8��(6oWoDb�S�b��$F6��I�l#��z~�K�����&1����ul�c���d?6�����lldc���X�F66���;ٛ���썐lr�\��썙l�d����:6��y�z�(E��:6oW�
��iٸ��U6��q���le�V��U6ُ��lފ޸��U6��q�M�d#-��m��ټo�ə�
���3�ټ��əlr&���79���lr&��Y3݆,�&��Q���l�'�ټ��q���
g�#�W�8����lgc8������M6f�<�7�7�mo�3���y*!Q�Q���lr/�٤\6)�M�e��F~6���m,h�����Fu6y���l�*�ټK}*�γysz�<�X�Ƃ6�Ro�g�:�ټK�q�ͻ������������dZN��%�}� xѩ������M�e�W�(�Ɣ6��1�M�e�N�F�6	��)mi#H���F~6γq�M�d#?�ٗ}oWor&�����y6γq�����s��N��Iȫlth�W�X�Ƃ6��S����&Ӳɫl,hcAڤS6����l|f�����lgc8���7oEo�g�:�٤\6)�M�e�i�dZ6	�M�e�<��Ωpd>ݼ��ɢl�(�,��pN�s���m��l�*����p6b����l4f�N����g6�%o�f#6�ټ�|*���9��M�d�*�h�&�����l\e�(!��FH6B�yx���$=6��1�ͻ�E٘��L6i���le�(E��C6��ɇl�!!��FH6��я����&C�y�w�*٤J6���l#���FQ6i�M�c��ؼ�q���l\e���&������l�{�H�FZ6I���lRi�H��U6��q�M�c#-i�H��=���l�e�*ٸ��U6��ne�(E�dH6o�n\�T�
���1�S�\�%H�l\e�*Wٸ�&����M�T�R�a�]��l�f#6��Fl6b����l�����U6��1���l��T�
�&H�l\e�*���������e���c�OiYږ�ұ�,���"��X.by���i�S�����~{����^Px�p]�ו����:�x��W\���3�gLϘ>�8��x=����3^1�?�띸����.����"�w�y����.�X������kl�؞�=c{�����^��eZ�������8<?�e�Y�������<��.�ɲ�,[����Sr�v������<c���9��l0����J��z�ɲ�,����J�ў�l0��l0��l0��� ��_��%?�ˏ���߻��������}�q_~ܗ��c�A�~D���������Gt��OG�Wr[�� �$����)l?�۝����������?�e���~�����g{�S��3z�� ��� �������lo?��������)��v�?%����?��?%��c�`�3��Sr]�uن�=g��ض�m����"2�+�s�f�gt���b�:��>ք[���?��?%.(�<��+�_��Q��S��$lCa�	��#lC�#�Lag
;S�X�������3�O:�N�`�Ӟ���&a7	�I�'¦6��)�M!l
��=���[���>Q� ��������?%���=���dw�]��}�l?�Ǉ���2�+�q?~܏���g���>�'�K���� �-��|��?��O�q?q��?����q?q�������ۂ���A>�����������p��?��O��������w��?|ǿ����×>Χ���×~��g��×>Χ����~����>�~��c��7�[�~Dӿ��W��6}
H?�����~��r��n��?���=������_�����l�B��<m
�B�������{��=�&�?ݹ���>�~5���N�I�mA�M�n����u\[�u�~m�>q��>q����:���s�~�p�&��qm�?��?���q��o����:����:�{��f��`�溙����N��5��;�k��6�k��~�p�9מs�9מs�9��q�u\�(�O�s�u\��nr}0�>\w��q}
�n��O��>��b<�����l���g�x��痖�n�����:���y~C�l0��l0�'����m�s���9χ�gz��gz��g�y��g�y��g�y�s�m�ن���g�yv�g7y��g�xnW���y���F�?��?%�O:�ǚ���A���ٙ������s7�lV�f���<�9ϧ��Y�m����Leg*{N�sʞS�����O�m�lCe�)~�nR�s�}N�s�S6����ݤ�&e7)�I�M�nRv����R��ܮ����u�_���|�)�t��J�7)L�`�'����;�����l0e7)[G��T>"�����ݤ���[�����H�֧�9�.m�i��6�n�ڧ�����m0��ݮ�ە��=��9��m0m�iL��iL�`��6�����m0��2�v��9��mC�SS��i�9��Lmgj;Sۙ�G���m����[��Y�ͪmVm�j�U��i�U��i�U��i�WۿڭOۿ����/�Z2�%C]2ԥ&������/�蒎�l��?�Q�]n���-��Ҝ�t������UK���d�K��d�K`��Ѭ��tiN��tiN��t��-���.��҉.���G7Y��%]������R������Вg��,5�R�.5�R�~�;K�	�L�=giN��t����|����ߒ�t	Lײ�,�Lk�d�k�gZ���g�Y-ېu-{�b��-e�Z<�M�E��Z�6�l0�Ғ��eϑ�.꒡�eZ�����R�.e�R�.e�Zl��Xu-6Hk�AZ�եL]����_�/�ֲ3-;Ӳ-�+Sr]vI뒴.I뒴��>g-{��uIZ�b�;��lCZإ�]۞���l�ж��j��vmې�vIm׶�j��v�c�<vJ�����h��v�h�v���]����]�f%�]R�%�]ۖ��]ۖ��Yit� w�o׶�m[ڶ�it׶�it�Fwm[�Fwit� wIm��vIm�vϴmi�إr]�6�mC�v	_��um�P؆��K���K������4��Ǯp�����d
ې<v�c�<via�v��D����]a��.��.��.�
�La�	��#�]a
�P�sn��'C������3�mH��Τ
^�WO+|�_�WO+ܒ�{��w�[����{W����]z�v9	� ��3�*x����w�Q�m�xI���5���į�Px	���g�����KN������Ka�������ؿ��ؿD�Kt<�?��5ڬ��K����I��t�S��9��б	���e��4�cg:v&��9��T2�ulV�f%�^ǇE}��G�c�:|�T��ؿ$�K2�$�S�i�C��3�x�襏^��v&��J�UڙT�KE��f�6+a��\��J~���+}X�Z/a�J�dZ�)yx�U�4��^i��Z/a�V/�RQ/��\��J2�$�K2���+���=G2��Rچ��KX��הּ�KX��6��^i�_���ۨ�a�A�_�k�n���S�X�T�K����uѵ)����� ��%�^��|^��%s^��u}��9���]����K����KӼ�w��R+��g[�������~�e�KӼ4�S������C/�� ?���O�[}�C/1�z�'���Sx�4�K����K��D�KN���KN���KN��߮h��vxi���� ??��O�vx=?������j��vxJ�ѿ��϶�x)���x)���x)���x	��Px��׳<;�vx	��Px	����@;<%na�G�������5�@t�ʿ�:�U6��!/��R��u��r�U�u/��r�%'^e7)[��xɉ�*xI����nR��ë�&r�U6���U��*��xi�W�y(M�'$�K������w��
^�%��gt���]���u���*xJ\c�B��n�@������� B�%����{��?�)�{��w�����{��w�v�lw�M�m
�ޥ�]J�%�]��n�e�K��4�K��4���<�v�lw	r� w	r��vIm��v����u��C��4�Sr]�	]���n]���N����{����)�^���n_���[ɻ5�[���[���S�4�m.��n��\mh+y��w+y�Q�ۨح��Jޭ�ݲ�)yA<�l�b���L���)yW�:r����[ɻ���e����-�ݲ�m.�6v�{��w�{��w+y���[�;%�Hg�F�nC`�lwkt��vKm��v���M|���)yF���[}���\ح���ۭ������>g��5�ۨ�mT�6vJަ`��ny��ny�6�uܺ�[��Sr�6��V�N�mXv �b��v��M�݂�-�݂ܭ���ۭ��R�m��6cvr� wr� w�o��v�o��vJ�A��X7gۙ4�[��;��-�ݦ�n����N���sԷS�!��6�v�j��v�c�<v�c��ۼ�m8�V�n��V�n��6�v�W����p�m����n��<���@�m���6+]�6vv�j������)�T�+��n��V�n�h� wr�I�[�;�*�*�ݲݭ��ݭѝK5�vkt�y�S�e��Tۭ��Jޭ�݂�)y'l0�ۭ��R�-�ݺڭ�ݺ�)�ې�v�j��v+f�A�[D�E�[D�E��8ܭ���벥�h��v����݆�n��6Gw��;%�h���n���n�u�Ѻ[���[}�շ[}�u�[W�u�S�FKm�i�۴ݭ����.�=� wr� wr� wr� wr� wr�a�[������Sr>�it���[���
�ǎ)�ݲ�m0��n���n�����[D��[���[������t�[�U�[�U�[��*�mV��n��6x�\�Y�۬୅��g�u�c�<v�c�ĝP�n��6x�W�Xu+S�)�[��M���v��߭L���n�6�w�I�tt�D�NtJ^�O:��n�v��tJ���՜N�{o��nꖡnꖡn��֜n��֜n��6�w�I�tt�;%.��q7�w�����|�m��V�N�E��s�\�� oS���u_��u�U��`�rݦ o�}��u�\����0�)�qF��-���n-���n-���n#�<v����[�:%Wog��nI딼F��1�[����ۘ�-V�7G���wBҺ%�Sb��nb
���n-��n��~6-���n�{�<v�ܻM������]���[}�շ[}���[j���[j����f�n��6�w+f��S�X~��ܮ�ɻE�Sr�	-�<�y��nst�bv�c���� 7"�]��v�j��po"��R�-����n�6�w�j��v�j��O�ܮHm��v�h��v��;%o7��n�{�ɽ[�����R�-��f�n3y���� ޭ����]v��V�n��V�N�E�`��ݺ�m&�.7"�n��<�mH������ht� wJ��6dL�.{�Fw�ɻ�[}��n�nj4�[��5�ۘ�mL�6�wӻ��[��e�[��e��0�-۝�����ܻ�#����m����n����n�|��w�}��w�������N�u�7��n��n��bv+f����)�.7"�ۭ���ۭ���ۭ��R�m�6w������)����[�)��14�!�AnrC���P߆�6t���]m�jCW���Ն�6D�!��oCW��)yFv!���Į#t���m�����Ն9����9���rCj��P̆<6�цB��0�6�a�m�c��	}"���#l��)qF#lC1��0�6D�a�m�jCW���Ն�6L�]m�jCW;%a7��Nɛ�F$Է���m���憡���Cs���P�7�����Cs���P�8��S�X�!���8�7�f�
Up���ݐ �8$���%ohtÄܐ�F74����n���ېچ�6���mC��)�.Sm��RmC��)�;�A�a�m�oC}F؆�6t�a�m�jR�0�6t�a�l�j�$ڐچ�6t����h��e�M�����k䫔)y�� Rېچ�6��!�m�h��ц�!�m(fC�����y���-l_#���-�<��D��)yx�+Z���N���T�azl�\C�*�P���5$�aTl�*�P���5L|_C���Я�X5L|�p�_C`��Я�X5��`��O�֡L��g�y(��$���LC`��}DR��uJ�Q���МN�kԉN�E�-0�5D�a�j(@C:%��A�r�r�)�aJk�rϐ{��sJ.�>aJ딼l��ttJ��O��4L|SZ��m�]Ǳ��W�xא���uJ.�c�k�W���)yx̱��\C�*�0�5��!|��K�3iaC�&��6��Sb]��)�.-l��ؐǆ6̅sa���P̆����_CD&�N�k�k��=�j�ؐچ��S��1M|��gt%�C`��)y��Fņ�7�����m�K��7Ľ!��m�j��lCi�چ�6������?!ېY�Sb���Ն�6t�a�k�jCW"��N���:��S����Nɛ���x�yp]~��������nH����5$�S�~�%�a��5��~}��>H]7Hf̆�S���1=vJ��g���2��е�htC�;%���p�0�6L��h��lC�����7Ľ��%o(yC�;O��fe��X��wJ^�_�<�
V�l7d�!�AnrC}��0�6�Os��P�N�3ڙ̾A�\�Os��N�u��L��o�}���07�����o�}��047�	p<�$����o�}C�z����7Ľ!�stC�z�0G7Ľ!�qo(y�8�)q���N�c��Q�F74���Anr�����N�ջ2�6d�!��n�vC���P߆�6Էa�m�}����A�a�mht��]�)(yC��� 7�ahnrC��憡�!ȝ���O�vC���l74�S�m�P߆�6Է!��oCW���Ն	�Sr�nD�!��mHm��OH};�?����	L���� 7�x� �0�wJ��}��a o�}�mC�0�wJ�	�L7����M��-�qȉCNr��v8�¡
3yC(B�
�P8T��
>��LG|T�G|T�G|��S��|�3�?���v�������LG|������mJ�UZڑ��\*-�(����(����(���hiGa|�ǘޣ0����	��{��G;|�����)y��Y���`uL�=:�cr��!��9���l}��x:���Q3y����G(|��S₴�S��^#��#>��#�=J�#�=��#�=��c��\��#�)�}����}����}����{���S�~�'$���ߣ�=Jޣ�=J�)yx65G�;%aS0���{�=�)yW��� ��9��c ����m�1�����*����i�Ǵ�c��\�mHN|��GN|��G(|�=B�
>��%�1G��{��l0�c �1�����G;|��G(|���Lޣ>��>��cr��6+��\��Ja|���0ߣ0>
�0>
��9
�>��#>B�c��1Z��{��G;|��Ǆ�#>&䞰�ȉ�P���P��{T�Sr�>"��CB�)ys|�	�>F���1G�(����(��䝰��{D�GN|��GN|�=&���Q��Q��Qr�����;%���9G�|D�Ga|L�=��cB��o���������{t�G�|t����c������B��1��t{L����wob��0�1��h�����j{d�G�|L�=F��i��G�|�=j�#:>��0>
�0>
�0��7�c��Q�����<�ߛwr�#'>&��p���h����GN|��GN|��G(|��G(|�=��#>B�#>B�#>F��u�v�h��9�G;<%�h�2mwJ�	;��GN|��G|T��L�c&�
��
O��v�dr�1��ȉ�����VB�#>����\�_򪂏���{�青��y� �#>�x�v����H��xJ��c& U�Q�u�������G;|���L�#'>r�#'>r�cL�\����cr�1�����ɽ���#`>�c��1����a�G�|���L�c���!�v�4�H��4�萏�������h��ɽǘޣ0��g�3ɉgG��Lr�#'>r�#'>��)y'��H����{T����#>B�#>B��lV��)yF;�*������G|�䝝�K�O��{��G(<%C;|���0�)�T���(����Gt<%��F�|t�G�|t�G�|t�Sr��4i��!��!������4�1�xJ.��'`>�c���4�0�1�xJ���(`>�#`>�#`>O�˖9��93�������#�>b�)�.�r�裏�����J���e�q�LO���,>b�#s>2�c�)[����t�#�>b�)���2���N|���t�|>��c��<�=�(�#�>��#`>�C����Ȝ���h���e�'�>�#`>�C�����w����G�|d�G�|4�S�~i������-M��4��&i�&O�ջ��&i�&i�&O�˶O�N|��G�|��G�|��G�|��Ǥ�V����ݐy�G�<%��n���#s>�c��4�����|��G�|��G�<%���XF$Oɥ�A2"9��S�]WJ����ԔLO�w]iD�<<��)yx�c��SE�*��G�L�SX�f+��:�֩�N�uj�Sk�Z��Z��ͩ�N�s*�Ӹ�C�?:f�����G�>:�[N�S2���)�.:f
�SE�*�TQ�?�c
�SX��9��:%�S���4�yJ���6%�.-�ש�Nau
��ı�iN�uj��4�4�9٩�N�u�ӜZ�4�yJ��/�S��F7�H{J�	;���iNs��Ӝ�|O�E�/L�w��Sݝ�4��;�ݩ��ʜ��)yA�!C��P�4�9u۩�N�v����"�9"�4�9E�)�N�v��Ӝ��mOɟ�]΀�\�/�v��S�=%.[�����m�n{J\��;��)�Nc�SʝR�r��;M�N)w��������m�1�9xNӜSʝ���m�n;u۩�N�v�S����Td�";٩�NEv*����f�mV�E�H;E�iXt�R��m�n;M������EO�˶3��|�a�)���m�t��S��E�,<e�)Ox)�FJ��;M���&�Ԁ�<�)�N�w)���4R:�)�N�w
�S��4x:M���K�O)�J�|O���s�S��9�Ԁ���)OYx��S>%�j�R�gجL�N�xO�J�4�zJ.�'ð��SO�J񔅧��S��O=�?�b�z�ԓ��|J��<uw�2�FJ�H;E�i�t����r�Y�i�t�2���|�)өOx
�S�FJ�<5�Sr����S��L�R<��N�x*ŧ�"�&�֡O��S)�J�T��,<��N#�S��𔅧,<�n�OxJ��d�Tw��;��S��ܙ��v��F7O�{/�NEv����4�9�֩�N�u�Ӝ�4��:�nNEv*����i�H;E�)�N����i��0�9�n����O�M���Tw��{J���a�s�S���4���|�*�4�Td�";��)�N�uʯSk�Z�V��:U�i����V��:��i2t
�SX���4,:��i~tʯ���4?:�Sr��!#��H�r���S��ݐ�;�)�N)w��&C��;M�Nuw����"|�Qw���i~t
�S��G��;��i2t��Sݝ��4:M������i�S���rO�k|H�)�75��Tw�_&W�75��4�9�|N3�S���Ԁ��;�)�Nuw��SݝR�r��;��)�N)wJ�SʝR�r�";M�NEv*��佷3)�S���6��NEv��"�i�";��)�N�u�=%�L*�4:�ճ��'$�N�tJ�S2����G���)�N�tJ�S2=%��.�|V��:U�S�4u<=%�_fQ�)�)�Na���8�����SX���V��:��N#����� i�Sk�O��:������h�Sk��G��:��)�N3�S=%~���S�J�S2���L���Sr�6��R� �׷��_�)ө�N�uʯS~����Z��:M�N�uʯS~=%�h�_��:��i�s
���)yF����)�Nau��SE���L�d:%�S�N��1?:��i2t��S2����4�i�)sN�sj�SӜf>���j���������S�=�<#��ʜ���}��W�|��`���
��Z����Z����Z����Z�J�����d�k��\�V��k�U>_��U>_c����*���yJ�	Z�C_1�C_1�COɥ�����k���L_1�U>_#��a�S�iiW�|����Keu��W}��Sr��k���G_S�����S���������"�r�S_���>������������䝰�k}��W}��W}M���諏���k ��L_}��G_}�C_1�5��꣯!�S��r�Z_��L_���<#����F]O�Eؿ���@쫵�fd_���Z_a��9O�u���*����
��Z�J��)�Wt|����)yx��4�ꐧ��M���m���
���yJ�	��!�W�|5�W�|5�W�|����+`�j�V�j�V�j�V�j�+M��L_S��4�J���������*����ʉ�)�ה�)y�ܮ<}u�Wa|���H�)qx��F9�5e�*���/y�`��O߰�=G�<%��細�H���ݮ<=%��֡C���+'�r�k��U_��U_��U_��o�:���r����
���+��?!��}Ž׀竾��2_���N�:~���WW;%����kN�U�N�3�5���|�[�������?|��+�Jޫ但2_����^��5��
r� ��o����o����o�9�W}{e��۫���۫��R�+����)�q,/�?�R�+��R�k(��^��N�k4��Jm����l�+Ƚ�۫����)yF��r���� �)yF����|�V��_wq�5���v�A�����)_qF� Jޫ䝒���='�9��+۝��w�䝒7�o;��W�{e�Jޫ�J�+۽��k��M��wJ���s�[��W�N���{��l
��+���k�� %�5"��{����|��W�{Ž��]��^����J���J�����j�b��c�<���|�C��7Ǎ���W1{�W1{�W1{�H�"�k��N�E�M���t|��s�^�[��<�}䫘���+��F$_y���^-�5��c�<vJ���a�U�^��]�^��^S��b���|E�S���h7"�_���^y��^y���^-���^��<��c��-��^I땴^I�\�,�_I땴^I�5Q�JZ�!�Ӿ<�}�`�k
�U�^�딸 ���^I땴^���^�ꔸFe�5���U��5�ѯ^��5�wJ.�nb
�<��yS�z��Sr�~ѨL���)ys܈�@�zM���)�.�&��+i���r�r���)�7"�_���uJ�nRv�rSv-�5Q��(<%�h*�&m���N�EHm���Jm����h���*f�b�*f�b��c�<��c�<��c���Lmjې��WD;%ogj�&�ث���_-���^-�5d��c���2|���D�kV�U�^��U�^��U�^��U�N�u�<����_-�5>�|���_ワ���j����j���Wj{��Ϭ�'�}��'�}� ?y��>y�3��<�|��6�O��ĪO�:%��c��N�3�M�~������O����O�����L�'V}b�'V}�ԧL}�ԧL}2�g&�3���P�uJ��ԤS����Os�4�Os��O`�t���ܧ}:�'
��gd���}��gB��N�b���O��O��T�O����O�9%W��]��$�O��$�S�� �'�|�g��[~܅�O�9%��F��=���}���O����O����O��L�}���r>Cs������}��>Cs�	�oنԤSr]�!�&Sr]<[=�u���Os��}2ԧ9}&�N�2!���ĪO����O���}b�'V}��)yF��X��P��5���O��d�O��d�Os�4���ܧ9}���9}�ӧ9�����eh�S�>e�S��m�3m����$�O��L۝��wϤr}F�N�Eؙ$��ݧr}*קr}*�g�F��i�O�L�}��'�}�>x�b�)f�i�Srn�t�OW�t�OD�D�OD���}��g����>]��>S��)�OW�t�S�}24�������}�٧�}�٧���d{��>�|�a�O}�ԷϘ�gL��>A��N�E����}f�>3y�lwJ�'Cx�i�O���}�)y�mi�b{��
��hL�3�wJ�	9�?9�3��ɉ��lV
�0~
�0���7nr�''����͐�g��&?i�&?s��Z�I��!�Sr]>���2��)����)��Q�O����O����S��&P���~��|~��|~2�g��\������Sr]>��;���S��G1�3w��;���Sb���)��C?s���yJ��.g��C?1�C���]N���Sr]n�,����.'���d�3��食>��t���Ϥ�g��S>���Ȝ���ɜ��������mj�)y�m
�?�\�}�(�i~��i��g�O(����)��I���M��O���Sb]��gD�SQ?��L?󐟊�������`��O���O�d�O��4��X�g��3���a<%��X�g��V?������������Q�Sr��!����Ok���OX���OX�L'~Z�g`�3��)�ߵ�]��"�)����O~�T�O2�����:�~��'�~��)����L��'�~�?���L?���G?��d�I��d�I��d��;��~�?��<�OM2�'s���r#�|���&����Y�O=%a�0Q�	�����D�g0�V?�3+����d���P�/w0?a�3+�i��d�食>��~*ꧢ~?a�3�i����i����i��)�Ok���S���s~� ?S��)����܈�����uO�r#"�~Z맵~Z�)�C��h���zJ^�mHk���OX��
~f?a�V�r�aV��G?}�+L�`T�OE=%M�h0�MT�OE�$�O2�$�O2��"~��g��SQ?��GO���IGE�T�OE=%�_�H��!�S�6��3d�2�~��)yF{�!�Ok���S�!a�3>�	���m0&
?a�SQ?���L?��3�	����	�������Z���������R+�)�S���)�.bJ��(�sɜK�\�)y,:@	��|�2�wJ��oDJ�\F����S�t�2�wJ��P���G����%�.�|�0�ٮ�.�+R��KE]*�RQ�d���%�.1t�[��2����%������L��{�<�C���K��Z��zJ.�L�[*�RQO�3����m��X����۞�0��%�.#K�]F������.u��\�����|���ݥ�.�}K�]��|����/��<#[�|�i���.uw��K�]Z��Z�Ѻ%�.�u�h�i�H�Dڥ�.�u��[��H���%�.��<<{�V���$�S�n���-��8��zJ\жu�[��L�����.u�[*�RQ��zJ.�nb�o	�KX]*�2��-�u�[Z�VO����v��>GX]&����Tԥ�.�tI�K2]��C��ϥ|.��<��1t��K=%��nh�2>��.�ui�Kk]Z��Z�ֺ�֥�.�u�;\Z�2w���%�.auE\*�)q'��%�.u��KE]*�RQO�u�U�e:q	�KX]��V�����Sr]vL��K�=%�jUd�I�e�q�t\��"���S�ܸ)�K~]��_���?.Evɯˤ�2ָT�%�����
�ˈ��Z�ֺ��'�.�uɯ���_&0O�3�\Z��Z�����KX]��2��T�S��W]���GO���`e.C�KE]���G�>��ѥ�.}t�K]�9O���_*�RQ���$�%�.�tI�˰�L�dzJ�B��a�eXt	�KX]��V��zJ�/7�Z��Z�)�%�.���<����͢.������Z����.���\�-�̢.��K~]���Z���e�ti�Kk]Z��Z�ֺL�.au�+��G���S��n��֥�.�u�����RQ�����.âK2=%����H��Z�ֺ�֥�.#����2���%�.�KE]*�RQ��zJ�/����%�.a��\�}BX]��V׵uh���R�ץ�.���X�����uݒ)�K�]�Z�H�٥Ȟ�K�K8�v�]b���%�.)��\��B��˨�Ҁ��֥/uw]7���|���Sr]�G��R��]�����Sr�nꞒ?4��x���%/Yx��K�]R�r׵��]��RwO�3�D�M��)�C��*�����ܥ'/#���)qs$�%1/�y��KO^�rO���T�Sr]6>�K�>%�jKS�����%/S��T��|J.&D�����evw)��ٿ�`/��K�^r����q�Sr�/{)�K�^r�z6>{^��R�����_ՙ^:�ҹ��}J.�.'j/Q���F���%j/�z��K�^��ҦO����I�^��2���%W/�z^
�2-�L/�{��K�^:�2S���e���\��O3_���̗f~J��]�f�4�e�y��KF?%�]N _j�R×��S��6+5|�����)y�_e�2��d�e>y�O^擗��%�/�}��KY_擗�~J��r��ۗ��S��2�2���e���<�-M _j�R×1�e�x3^2��ї��e�x�<>%�eK3������/e}Y>%a��O�uٿ�:/I~I�K�_��)�.��p���%�/�~�>%o��;�ԧ��m����se�z9*P�
��Sr��ն�:cP�������A9c0%��ӯ3e"z;P��mHz;c��L�E����Ǯ���6$�;h�ڱ�v�;hg�{�v��\o���vƠ�`og��vƠ�`o�ڹ�v.��mnz;�&������o����L�E����ag5%oۨ�������m�z��ަ����-�oy��<#;�^6-�����������-�o��[��Ʋ�J�U���oc٧�5��j-��']�f�ٚ���(���ؒ����m�{���L�u��jGڹ�v�oo�����6���h��!�v��m{�����6p����o����6p�h� �!�v�Io� Z�ߊ�V��Q�m�z;���C m���\�mȹ�V����mnz����C ���e��q.�h� �!�6p}�t=��3ا�ͱ�8*Ў
L�E�Ar��(h�ۧ��_���c��A��ގ�m{��ގ�3mnz;P���s�\@;��C �@;�����mnz��[��F��Q��@;��C m�z;��w�8�Q�vT�h� �����h��۹�)y'l��C Sr]�G�ڹ�v.�h� �!�v�Mjo���R����6Q�ڈ�v���xog��v�`J.�Vk|;v0%�����mR��\����v�o��������(�V����-�oy���(�6J�h� �!�v�h���<�����s�\@��>%a2]��h���6��(h
ځ�v��hGڹ�V��!��oy����������!��o�}��[F�擷��-�o}k��|�ѷ�孬oe}�b����ѷ�~J,BY���ؾ��m�y��[l�b�Nې��S�&�oI~K�[��f��J�U�m�y�u>%��J��Z���O�Eؙ��mHz�������S�>R��*mV�Q��@;0%�e�r.��h��O���C �@;�f�O�����N�C m�z��ފ�V���MWo� �!�v��-�o��[�ߊ����J�U���o��[����V�JJ.�fe�z��[Fߚ��̷@��-�o�|�[ ߆���u�-jos�[��榷��m�y�ܧ��&&����-�o�|��)�.��譬o}��ې�Vַ������o���\��IF�2��ѷ��e�mx��X�������o��[l�b�۷ؾ����o#�[l���Vַ��Sr�$���o�}��[l���Vַ������o}��[F?%a�3�5�o�|���2��̷f�5�m�{��[3ߚ�)yx{�@���S�m|�.'����â��𭆟�g��Ϗ&�O�u*�&�O��*ߒ���	��o��[����O��]-����so�{��[�>%/�n�Momzk�[��湷6���-Doc��X����\��=���:o�y��[u�󖘷���x���)H�[b�z�֓����so�yK�ۈ�6Ͻ�somzk�[��F���`������
�6�E�-jomzk�ۈ�6���-Wo�z�է�lC
�V�����m\|+�[��r�֦�6���S��Mo!z�[�ު�V���U�:o�y��[uު�Oɥ�j%�S�>?�M���6쾅�-Do!z��F�O�g�6�+-K�RX:�.��^��<�o/�Ji�)�v���~[ڔ~7H_�3�����]��L_ɥ�v����;�W�~�Ӿ�K�mC_���mC_��m0S�m0_���&_�����)��������W�`J�ۨ�����W�~�6���?�_�3�~ܿ���g�w������%Έ�����W�X~���_��U"޿�J��w���	!ſ�g���|%/�w��\����+�.�	,|J�_�|%a���%����+��		�_�;���J�ў�'�J���+����m0H��R���J�U{��+y������~ʦd7YvX�W����J��6�'�J\#��_��o;��+�z��Wb]��%��F<���F���}N�J^�;��W�mi���R�r��E��Wrn�ș�J.��+�r���rd�O���+yF���_�3�~k�������J�h��|J�/X�W��A"g�+yAn���_���!ſ���3�¿��J�������|%�egBw%n4A�_�Eؿ��J�{�Wr]�4�W�Nج0�_�3ڬ��_�3ڙ��_�;ag�r%��.���\�->%�,�+�z7n����m|���ܸ�?%wiP��ܒA���!��+y�l|��%�e/D�%���JS�)�����R��g�e{<�G �W��@��ĝ �%���+q٨��R����+y,[,�+ys|2<n�`�_�3�kB��W�!�ῒg�!ſ�gtE���|�Cw%��<���5��"�}Jv&�ۿ���3�d��)نP�_�;aB�%a7�%�[2<�W���_��&��+���W�v��Wrv�W�n���R�+y��0�_�E��"��+y��/R߿���3�¿���Y!ſ�?m�A�S�Y!ſ�벥a��d�|%o���%/��D��W�Xv&�W�����%���P�����FA̿��wD�J��Ol�Wr�� ����+qF��W��$�%�	�S�� ��\�Ϣ���l����"�ѿ�g����<�����<���>%{!��+�T<q�_ɟ��>%)I}�J����s����/Π�_�{o/Ĺ%o��������m|D�%o�-���\�-�����mC���/��1u��X��_�E ѿ��%�j��%~B@���Rmi@����_x��lVx��5ڿ�s��=O��<��X�����F�d����+y,�3"x�+yx�_���m0���ݒ=�x�+�.�dx��"�L�΄'�J.�sg�'�J�΄'�J�)�����������(����� ק�>�����"�� ſ�)��<�Os��%�݄����&�v�D���]u�1�J.���_�E؆HD�J����r��M�J�hmV��)٬�R�J.�o�\�J.��j�J��6�`�J�;�	���<�=����տw���X�|J6+��W�Q�_�3ڬ�R�J��;aKæ%~�D�%�n�����5��P�_�k���-u��\�͊`��R�9H���}���%�j���%�h�Aw%o��mO��A��W�>��)���8���>����M�n�t�K��t�K��tۋL����%�^����Z��EZ�W�����uL���jJ.�/ŗx|F��\*=g�ɗ�|�ɗx|�Ǘx|�ǧ�"x(���`g�H1�J.�f�T�KO�H1�J�=Ӕ<#���M͔<�i�Ǘx|�Ǘx|��a�_��VKb���K<��=G<���S��,�J\6��_��Y>%vCK���'�J.�M_��)�㐫O�u���ꋬ���_
�%W_���M_�%��j�gZr�E��Wr<�-�����Eج��K�>%�Ŗl����_�3ڿ��K���S��r:��s_:��`_d�%oK#�|J�4��ҹ/�R�/����/"˧d�!��+�̶�H̗�|I̗�|�Ǘx|)�1�_�k�)h��|i��|	���{J^�@��K�ߋL��pS�y([Č%a� S�+�[�R|)���_��eS y|Jn���K�4�� ���m
��E��W����¿gT�/��R�/��
{N�s�K�����Dʽ��K�=%���Dʽ���J.�6Dv�W�m0R�%�^���^���^��%�^��%�^Dp%�hRdO�˶爴���m�C��t�K��H�_-E��_/a�V/���LO�����:T�K���K��ы��)�M��K����������C��W��&Dp%�e�!��+y�6E�Rd/E��_/��V/a�V������5�!\�+yx���zɯ��z	���z��\����\�����R�9�~%�Ï�z���\�͊�)��9�/��<"��"��+�za�"��+�Ta�V/a��\�[R�����Yi���_�Eؿ��KX����J��6��!���Z/��"��+�.�>��%�^��%�^dw%�e��_/�����r���G�����=궗n{J.�^H��W��B������	���{	���{	���{����zi���z���X��z���X��z	���z	���z���\���q�L/���L/����gtKv�	���z	���"l|Z륵^Z륵^Z륢^D�%aK�LOɛ��MX��ՋL��Ǻ�9v9���\�]N~�#�J�8��][��_�˶�����_�3ڬDڋ���ݥ���<�]� ��e�͖�{I���{ ��8�H{��׳궗n{���H{����R����\�[EĿ��c>;�n{���<�� �)����Kݽ��J�	;ӳ3=;��_�c�:��Kk���KX���KX���S��ĭ��zi���|�Z�g�!��+y��9"�^dw%��^dw%A��W�樻q�S������{I����&��%垒w�-��_�u�`�gѲ��,|�)��\�[2��"S|Jv&���<��I�=%Wo�Rw/u�*�L���^$�%�6Jݽ��K���KE�T�KE��}N�s��KX���KX�Tԋ��čV/r���"�+�Tr��d�Qd/E�Rd/E�Rd/E�Rd/�¿�����"{ �i�_�3�Mt�K��t��;Z-��.o�=Gݽ�݋L�����K��J��@Y�������ٙ��$_��_�~%����_�_��%�^$|%o��P�H��J����x��x�䝠�n���o����Ɣ�rۄ�m���q��<#��˓��{�R|+ŷR|k��|���{����{����[ݽ��[��u��h�m4��rq#��l�>�l��?����n��ߺ�oXגg�o����[ݽ����%A�ق�-�ނ�o�ɒ?G�7�cɥ��sظm=�֓o=��o���o���)����oS̷�|�ɷx|+ŷR|��?�h�˶�·,|l�����fϴ�ݟp��-��-��F�o)��ro)����,�qx�*��[�,����m��րo�րo��VwߥX�GY���Oז��c�ɷx|�Ƿ��[<��?�Ɵo�Ϸ��[u��:���Zb�헒-ͬ�-W����M�B�m���?K�N��[��6��O�u�,�E�[���[��M1ߢ�-jߦ�O���O����[����S�'dU�o5���o��6$}��!�[Ծ��o��6O�ې�mH���BQ��<��J�>%���I���?ߢ�-jߢ�-W����o�ͷ��[�>%a�2�|�᷉�[ ����D�-��Ɵo���\��4���o���o���O�;��NF�I���-��2�-��2�-��2�-���o�6�|�跌~J�	[Z�Ҕ�S����!�[?%0|F6$}�������f�oI�6�|l>%�ӯp�u>%�e��o-���o���o���oŞ�5�r��-��*�������������I�$K�$��U���r�v&��V�o�ϷJ����5ڙI���-��Ɵo�ϷJ���J���JJ^�mH����[��U�[�?%�e��oI������3ڬT����mn�67}������mn�V�o��V�o��V�o�Է�J�]�Q�[˿��[�����(��埒�m/��oCҷ�J�f���*�)y��[����[��%�Srv9���o���o���o���o3ط��[����[���e�Z����Z�m����oy���oy���oy�6�}��\߆�o���oCҷp�����[˿��-��6�|K���S�@��U�[��U�[���?���)y��r��-����m��6�|��)�[��%��`�)y'|���oI���O��ۙ��S��ؙ��[Y��:���������O�跌~��)�S���[3�5�[3��:���m��6�|�b��[ ��[���[���[���[�>%/۞�� �ܷ�����`���裛��Sr�6�ȷa�[�>%��n��'�[ ��}��m����o���8�7�}��~�u�6�b�����֡����m��V�o����oQ��oQ��oQ��O���}Y���|�)���t�[ԾE����`�
��`�
��`�
��`�
�m��V�o�V�o��6�|+طY�۬�s�����ج�����m���O�u��Q�o�Ϸ~�u���[��:��m��6�|��䝰���󭿟��r#���7ǯ��'�����������������������m��V�o��\�]NY���[F�e�[F?%�e�S�o�η�~�跌~�跌~�@~�@~�@~J���'�ߚ�m���\�Os��m��o��6�}���%�[����[��`�b�m���o��6�}���[l���[3��[ ��[ ��`5|��C�O��������O(���BY��)�މۇ�>��aR{��Cl���̇f>�M�����Q�!��}(��hV!���w�fF���>��a�z��䝠3�$?\��� 4�)�T�U�Ʋ�C �����b/7%�EK�¹�p.`J�����s�\@8����O�3�1C�������?������C���0�=����-h�C���0>��a|��C�������?��Sr�ZS����P���?�x��C����I�S�l���P���?o� �!�P���?��Sr]�Gy����6>�(���5�������?��!�y��C��Ň�?̆���C������9�����X�C �@���ďC��ʇ�?����-h�C����p?L��~�F��P�JJ^��B�}��C��ۇ�>����e}� 2�0>̆e}�fÇ�>��a���\���P��߇q��}��C�����>��!��}��CF2��ч�>�}h���QF��0g~J��˶���DY��Pև�>����e}(�CY���̇f>4�S�n��a�|h�C3��0z>�S��ۿ4�!��|=j�0�>����C��0�>D�`��C���0�~~	�F���Xױ���Cj���O�E���Sr�4�|��߇�>̿e}(�CY��Pև�>d�!�}��CF���qgu�YwVǝ�$?$�a�~��C���p?�������\��Q�Z�0�?�����~�Cb�0%?�����}���,���������C���08?��~���������ר��}������߇�>��I~H�#m�&�p?��!��~H���P釉�a$~(�C �0�>4��|h�C�:�����`{��C���Г��<��a6���]��g#�"� ���������!D�$D!z� &ȇ	�`C��� ��)y�� �ч�}J�ѭ�6=��a�|���P����\=��!W�z��C�B�0A>L��z��C�&ȇ	�`�z�է��ݮ(��l����=�a\�����3]ېA�!jQ{��C�������a�{�湇�=D�`{<{�I�aR��<�F�:�й��=t�Sr]v&��C�湇y�a����8�7�f�lVF���|h�C3�)�;�@>�a���\�$e}(�CY?%��6J �PÇ��a�|��P�0T>d�a�|(�CY��0g>��S��h�z�/�d�����>���}����O�2.>����e}b�ۇ�>��!�S�CF��0�=4����\��KF?%B�4e}(�CY��Pև��!��}�F��0�>$�af}H����P釙�!�I~H�C?%���d�)ys���([m�W������C�f�O�E�m����@8��s���(�C��������!���C�������?Ώ�!;�C a�~8�C ���\�;QG�Q�pT ���pz ����pz ���K����
���@8*��s�@8��C S�Z�¹�p. �s����"��v_���p� ������0�?�D����p8!�;0�J��8N"L���S�=�q��8cp�18�L���cǱ����q��8vp��j��R�����p�1���?%�J�=N5G�#��)�.���G{<�+�p�W8�+���8�0G�#Ƿ
��#����q^����$���������S����8vp�18
��ٜ
��8�g�3���@��}��� �Ǘg�3����q��8P0%�j{t��8cp(8
��؉N�[h��� ǁ��@�q�`J^�]���[�c����q��8*p�8���sǹ���Q�3��C �!��lV�Lɟ��iٙ���7G���Q���qT�8*p�8���sSr]�4_p�8N� �C Sb� ����9ۖ���qT`J��f���qz�8=p8�
L�3��vz�8=0%o��ʁ��@��� �����cǱ�)�.�r���r��$�q���?�?��5�;%��C�qaJ^�����p\ϵ�7�p�j8N5��Sǩ�����ǩ�)y'��9�pN8���r�)q,���	��� ��
���$�	�9��g�3����q.�8p8���� ������O��fJ�q�������c��Q�y�1�������w�����!���q�80%�nȹ�cp��\���cp�18���18���cǱ����q��8vp��?����1J,�!���?��������90%ar�8p8� �C G�T�G���Gl��S�چ��GY?%agR�O�E�]����1K�H������c$�Q���Q�O�E�҄�G���Sr��4�����1K���pJ��Τ�?�������I���I���I�������������$�H����������)yF7[�O3�N�P��4��C Ә<�]�!���?��cJ�1%�8p��?�
#����c��1��8*p�?����-�u80%�e71�~J�ޭO�`(8������d����qz�8=p�8N���ǔ��\�q.����?F�
�����cJ�q��8vp;8�#�cS�c��^����I��$�q�8�pL�?'���	�I����q�`J�����I�cp�q8�8�0�?����(G�#�\��T�q��8�0%Wo_����}8������9q�8�CL��e�vh���8M�g�v���r���qBbv�ކl��q�bJ.��=:mq��8�VG+�/8�Q�p�8M�&��8M�&�o8�Q�(�s�q��8�q�8�pa8�0G��
�7G��
�y�c����������ǩ���q��8�pN8'�p�W�����8�pa8�0G�#�W�����r��8�p�}8�h������q8�8�0%�j�0�J�͖�	�@��p�q��8vp�18G���Q���qT�8*p8����������?��c��Q���Q�C��C �!���?�>�!���q�80%�nȹ��\��\���!����s�7�p�8� ���ǹ�c��q.�8p�?��#�?��cT�����O�k��/-���-������e�Q�e�Q��������Q�Gl����#�������������(돲�(돲�(돲��菌�h�f~J�f��?j���?��5�Q��?������̧��)�O}՟2��ѧ�>�)����`�����\=M�O!z
��x�Ԧ���i�~*�S��B���=��)DO��Su��4�>ͿO�y��B�4?��iJ~���
�T���=�`OS�S�>%�EgJ��S�:�Թ�Y�)}O�{��S�:�)���6=��MO��Su�&ۧ=��)DO��S����T����i�}
ѧ�eۿ���<%�'�e�Zl���٬��J��&ۧ��i�}��S����)�.�A����3i�S����Ԧ����MOmzj�S����Ԧ�6=��)DO3�S�����T���<��O=y��SO��̧�<��S���Srv&�x�F�������)�?!=y��S<>%a2�>%�)1O�y��SO���4�>��'Oc�S)�J�4�~J��4�>��'O=y��S>%/���Ԁ�<5�Srv&xj����|��;M�Ox
�3lԧ�;���	��Ӝ�4T~JH��̧,<e�Ox*�&ȧ�;��Sr~D�s�p?!�N)wJ�ӈ�4�=�sO�w
�S�R�)�qx��'�ݩ��g[���Tw��;��i�{�����m�n;u�)�N�v��S��"�i�y�i�{�ӈ�4�=�xO�w
�SݝR�rO�3�Mt۩�N�v������O�Ӥ�4�=��Iݝ��4p=��)�Ns�SݝR�47=��inz��S�=%�ѯe�ݩ�N��S������;��)�N�v�S��"�i��:�mH~�Z��ZO�k���O:��_��:��)������m(mC���;��)�N)wJ�S��"�iOɛcg2$=E�)�N�vj����3��I��"�4�=٩�Nc�Sk=%hv&��\�&� ˞Z�4�=��ix{*���R�L��4�=u�Sr�v&#�ӈ�|��;�Srn���)�N��Sݝ��rO��m�H;�i�{�瞊�_��:��)���䳕�:o��g���:U�i�{���Z��Z��:�֩�����Y	��<�V��zJ����:U�)�N�sʜS�2�9��yJ^�mH朚�4�=5ͩiNMsj�SӜ�4�=5�)`���4��yJ�˸�T>�q�i\|��S����T>��9��)sN�s*���4A>M�O���"셆ʧ>:����hK3�=�)`N�\�{&��S��f���9�i��<�{&��\��I����T>��y�L.��41tޞb�4�=��)�NMs��S�<%�%`Ns��S�<�G.H��j�4�=��i�z�S��:����):N�S����4�<M1OS�St�����8�i�x�������8E�):N�q��St�����8M���j�!Oɥ�]�&��8E�):N�q�O�:�4�<��)MNirY>%Vo�y
�S��j�T+�Z9M1O�r�b��4�<�'Os
�S����&�49u�i�x�� �4@<��i4x��0��9�)`Ns�Ӵ�4<̩VN�r��Ӵ�0Oɛ㞩�3ɜS�<%�j�U>��9��Sr]�Z1t��S�b�)yx�g2-<MO}��<�S2���4S<Uԩ��*ꫢ�*ꫢ���O�J����)~����+����k��5f�
�����L񫵾�_ħ�"�W�}��f�_���mO�u��R�+�R�k��\*�j���j���j����<~���)�v�W)~��W)~��W)~��W~5�W�=%A����+������_���rO�3Ґ���W�}��W�}����+���V�l�f�_�ί���|�+�����+��&�_�ՀO�3�De�W~5����k����_Y�5y�*ůR|J�	ۣ���ɯ,��¯)�W~e�W~5�W~M1���_u�Uw_�ȧ�ظ])��m_3ů��*�������k��i�mi_��i_s��n��~����+�R�)�.�_��+�R�+�F�O�;a7|_��Uw_��i_��5�궯n�궯n{J�	�Q�_s���{J�n"�R�k4�UwO�E��1��~����+�R�kv��nW�{S��n���vo�ݛl�&���k��Uw_㼧�5j���j����W~���~_��5��ǧ�Oȴ�+1��+1��K�Y3~%�Sr]>,�Χ���R��v9#˯��7���K�~E�S��/�ͯ��W�:��+���+���K�aѐ�����k"�5��诌��诌���~��WY��WF�M��+����_5���_#˯�������}J,��1�7��U�_5�չO�k4�����"l|j�����gt������+}��ǲ3�ڧ���L:�)y��Lj�+}���k���\�_*)د��*د���O~�'��O��)(دa�W�~E�W�~�ט�k��չ_cƯ��J߯��W�~��Sr]��t�&}�gT�_��M{���J߯���O~E�W�~E�Sr�!#˯��J߯��Y~�,��L3���|�)yF��,������j�kd�U�_5�U�_#˯����򫙿��_�ȯ��
�a�W35�W �W �W ��`�+����r�6>���_5�U�_ѯ���D�)�._�Ī��������7�*�!��D�+��&�_��5�J����u~�:���+ɿ��+ɿ��k����_�ίY�W���W��W��Wl��Wl����+����{�_��+��&�_e�5S�*믲�*�i�WY��״𫬟����)~��WY��WY��WYM�b�����������)qF�����n�t����+j���k��5��J߯���ܯ��W�~��Sr]�C��f��}��2�+��j�k���O�[��h�+����+����w������m��W35�W35�Sr��gR�Oɛc��_cƯ���L�k��5@|:-�������������������_I���O�E�A*[ZٿʇE-���9v9�ɯ��Sr�/��s�|�)y�>:*p�����b>%���3����u��:PpM1��w���@�����:��g�:vp;��\g���Q���uT�:*p�'��\��U�_��U�_��U�_��U�_�ǯ��j����W�U�W���-����=�L�ҿ*��ҿ�_��5@�j��p�
���R�LZ�����+ܿ��+ܿ��+ܿ&�_3ů$�J����������å�M��WY��WF?�?�5چd�WF�2�+��2������)y��9�'��'��g���~��3S��)�d�OF�d�OF�d�OF�4����R�Y=���?S̟��)럲�i�f�i���O3���O��t�O��t�O�����|�'Wr�'Wr�'Wr�'W��gd�3���՟\�Y��O��L1���`
�gd��?Q�3��Y�t�O��D�O��D�O�>%��f�ڟ��)؟�}J,���`
�g���?S̟���ڟ���ڧ��L�-ٔ<���`�s:��s��'j���`
��`���b��LD:��s&�?����O�E�u�O��LD�������6��ǲYi�f�i��l0�c>��O���M��`������'��g����?����?�ϧ���n�LD�f����'���'�&�?��3����f�i�@~J��6$��?��3��m;�v�&�2�'�2�'���7ǽ����>%a�27�)��5ڿd��D���Ɵ?���?�ϟ��O��6$��'��'��'��'�j��s��gH��?sӟ���ڟ����t�O��D�Srv!�S�?����?��S�?��3J��ǟR�)şR|J����iJ������ɟx��ǟ,�����O)>%�>�X�g,�S�?���\�����O��oB��:f�?!��8�6}J\�6�iӟ6�iӟ��O����O�>%/�ݐ}J�ѯ����<��`����>%��I���s�?5�S�?5���?����?Sߟ����t����g������c{��?����?����?���f�	����~J��wl|�'}ǖ����g�S�?5�S�?5�3.����O ��j��sF�?��ӹ?���?Q�3��)؟��)؟��)؟�ψ��sr�gR�ӦO������O���O���O���O���S��������ܟ���t�O���O���xr�'Wr�g��S�?�S�?�S�?�S�?��3�)؟�}J��l�g6�ӹ?Q��?�S�?�3�]����O����O����O����O����O�����P�g��S�?C埨��՟��O����Sr~�%j��?4{���O���&�O�E����g�^�@�	�i�O ��O ����e�@�	�@�	�@�	��π�����K�c�蟌��蟌��Y���OY������'��?��s_hf�3����O����O���Ϝ�'�b�)�z���������F���Ol���Sr6�g5��=;���i��p�	��p����J��l���S�G-���?���?��J����$�I��������d�g����?I���?I��X���)럲�)럌��l?%��^Nl?%�e�R�?e�S�?�����C����ퟹ�O���O���O�L�������'���gt{����w§_��������@���b�)���������������@�g��3�J�8|�5�����$�S�6>���p�	��p�	��J����J�1�0��i���"���\�g���?���������O�����g.�S�?��S�?y���?y���?-��?��S�?��S�?��3�����������'���?��pJ������)�C����D�����'���g����?����?c�1�%�/I~I�K�?�ߥN�w]%�/��K�_��R����/�|i�K _�2z~����nR��R֗��L�/��ˈ�2�}J�Cv0%�/�{I�K�^:�2���`/�{��K�^:�ҹ�νt�S�ׄ�S湗���/�{��^j�R�O�uѬJ _j�)�.�>%�����3��^������}J�Q�^�����y�%}��P�^��)�;��%�����	�K _�2⽤�s/Q{�ڧ��V:�2⽤�%}/�{I�K�^��2���e|	���Y�@��%��e�3A�d�%�/}i�K3?%�-m�������-[�$�$�ef���_v9�~�3_��R×��D�e\|_:�ҹ����S���ˈ����\���e�{��K�^r����y�`/{)ا�l0
�R��6�L}/�z��� �2����S�m
ۦ W/�zm��vc6|)�K�^�����/S�K�^������D�S��M�����%}��AJ�^f×A�/S�K _���y�%j/��K�^Ʋ���Lj/c������쥆/�K_���Q�%�/�|��K�>%�h됾�νt�s/�{��ː�2$���%}/�{I�K�^:�ҹ�νD�`/{)���2��t�s/�{��K�>%�e{I�K�>%n����I�^:�2����%}/����>���K�^���������O_j�2�}J�/����%}/�{I�K�^��)��_�����s/�{��K�^湗\���S�v��WO�.g|I�K�^����Oɥ���e6|��K�^������앶4S�K�>%/j/S�K�^F���}J\��牢/��K�^��W�M��!W/�z��^f���%j�����>%��.M _�R�Wچ��%}/�{��+ݥ�ڧ��L
�R�����e{)����R���%j/Q{��K�^��J�_r����\�\/mzi��t�����\/!z	�ː�2$���S��6�z��K�^��Ҧ�6�T�:/�yI�Kb^�2$�I/�y��Ku^��R���$�%1/=y��K<^����x���%/Yx�^�𒅗,�ߥ�.�v)�K�]���Z�����%�.��K=%����g0żT��|RQ���e>yI����RQ���T�%������.�.�tI�K2]��C����Srn��%����]=%��Ï>���������`��G�>���e�y�u^*�z�M��e�y	���"�9Z��Z�Y祵.au	���ܮ^Ɵ����?/��K�]��2���%�.�u�u^��)�.�H��e�y��K�=�?�ͱ=��K�=%�j�i�H��%�.�����Rd���6/�u����L���S�N��,/u��KE]*�RQ���T�e�yl^������ե�.��KX]��V�d��:/����K�K2]��2뼔�e���\�F�\��R+�4���S�3^��)yF?��0OɻjS�9�1�e���<�M��3�K]�I]b�R>���eyF^���a�%���g�F�ARQOɥ�A�Z�ֺ��%�.au	�KX]f��ֺ�?/�uɯK~]Ɵ�ֺ�֭����[X���6���m�y����Z���m����l)���_����׭�n��[X=%���c���"�M1oS���)y��n���m�y�[��Ɵ���ox޲�ր���-o�[)�J񖅷�5�ox�[��f��໥�m�y��[��f�O�ó�j�v�b޺��m�n�uۭ۞�Xl�ڬ�|���-�nuw��[��R�r�����-�n)wK�[��f��Y�-�n��[���(oxl޲𖅷���-�n)wK�{�Ҥ�-�n�v�[�=�f��L��i�Y�-�n�v��[����V��zJ��δ�L&����m�y�Ɵ���-�n�����6�|J��Τ�n��[�݂�6�|J�	�ٚ��m�R����-o����򖅷,�e�S����h�Y	����|��#o�w�[�݂�|O�k���{�s4�ou����6#˧���_�s4�S�lC�6�mCJ�6����-oYx��[��R�r�����-�n�w�����6���?oYx��[޲𖅷,�e�-��+�V�O�3چ��-o��[O�a�2]���'o�x��J�V��R���S��|��J�V��R�Io�x+��D�)yF�4�oxk�[�=%/�6�nH�݂�|�Y�o�w�����O�ox޲�O���,�e�-oYx���J�67���o�xk�[>%a�3J�e�m"��<�]N޲𖅷,�5�mHz��[�&��q��o���`�V�����-�n)wK�[�ݺ�6�|J^�]N�=%��.���Oɛc/|����md���Fx�[�=%a�ҀO�uٿd�m"z���D�6���m"z���&����:o�y�󖘷ļ��'o=y��[O�z�6]��Ro��[<���67���S�N��LWo�է��q�g�z��[uު�67���mnzK�[b��)yF��%�mnz���B������m�z��r����\��M��R����MWoQ{_��ν\o�[�j�)�T7�j�V÷���mx{�[�&�O�u�D�-�o�|���V÷���-}o����Ѷ�������o5���Ѻ	�O�u���u�(�o3���۷쭬o��[Y�F��Q�m�z_ۣ����m"zޒ�6��%�-�o�Χĺ��P����������o�~��[��f��Y�-ɟ��w�f�y���`�~6I~K�[�ߒ�6��U�S�F�qS�)�-�o�~l>%a�R����o�~��[�ߒ���ؾ��mdy+���}��ѷ��-�o#�[Y���6��������۷������o}k�[3ߚ�ȷ)歙oS�[ ��6ż5�-�o5|�����)yx�P�ϑ������S��L�6��#oc�[ ��6y�5�m�x��[F߆��@��-�o�|��:�ֹ�νo�{���h�6�u�so��[�ަ�O��@��-�o�| ޚ�6S|J,՘�n��1�S��<ޒ���O�E��T�m>���9�4y��[����V�J�%�-�oI~K����9�mVm��򷖿����oS�[�?%�h�R�a�-�o�~�[�����J�U���o�~��۬��߷ؾ����o�|�O�0����Ja)-]K��o��J��|�?�U�����%/��i�+K��w��\��3�Wr]���+������"~�g��o��J��}%/�wg��������<�og�J��w����8������Wr���+��ߖ���q�>N����+�����W��T�J^�o��J^����+������\�o��J^����+���.��\����+q'��.�+��e/�%���J.�^��J.�w����_`����Z�U׿��������������\���l�(���O���ˎ	��J���~�E���ގ����M�X��䝰�����\�}�?��M�Wr]��e�$J}Jv���/�J��7�_����~%B�U2ؿ�벯.�*�_�{���ܔl�����m�|%a_e�+qF���li(����_�����_(���"~�2�������d��n�-m�Ұ�_ɥ����J.�M ��+�[��+yF���+y���J�	�׶1�\��B���Ku�����%M�_��%oKcz�+yٿ���+yF�_�kt�Ȍ�Wr�/���wi����������J����<������F�	p�+��_�0%�	J�+���%o� ��+y���}%a��O�>A��Wr�,�Wr]�x�Wr��	��W���s�J��ց��J.­O�:��_�û���%o�}���8#J�+qF��W� �_�����J�B����Ԡ�d뀾%��F������n}�J.�+����?�J.�]��+�T;���ܿ�gt�>"����\��Hd�%Bv ��W�v ��W�N�' �_�u��@�%�e7!7�+�.�>������ĺҞ��J,�t�)ن�R�J��6��J.��tτ��J��m��_�u���Oɝ��_�c�� �_�rτ��J�2ٿ��_�3�A��%/�f�6+��W��X^�--mi�����mV�%o��%�;��3�ڿ�?!;\�+y�mC@���e�����ll�Wb@��ĝ �%�eg¦%�j�"�}J�! �Wr�! �Wr�!�ڿ���΄M�J.��W��Os$�%o�¦�?��eۿ�e�J.�f�M��7��Wr��4����Ld�%��<��� �׵A̿���fb��\�-����e��ѿ��rgE6�W⌨���A�%A��Wr]�4l�W�;+��dK{��g�B�%a�"��+y'�_��%o��Y�ῒK��=wi��O�^H��Wr��g/$��+yx߳���g�N�1���J�8|�}>�b濒�r��J�Ѿ���J^�}3��<�F���8��h�D�%�l��\�M����R��_����l���)�	,;&��_����%a���O�&Jf�W�'D��W���Dɬ�����<��4���m|(����(���"�����?!�(��+y�l|��)�U,�c���_��vCI$�Wr]>##���벉�M�!���Rm���Q�����OɎI��W�Xv9x�W�������_�k�%ܟ�������W����%��ƭݸ�迒w�6�>�����\��4��Wrv&H�Wr�!H�W�N�%C�%o�!�+y�n�0�_��� ����~���J.;�_ɛcS��%����+��u ����_���,����O�w�K��$�K�����J������J���ג�/-���/��R�/I�"��+y'�Y-���/e���/꿒K��,�"�~J�s��~�藌~i��}Iߗ�}��A�_��ӆA�_ɥ҆A�_�_&�&K����l����LK ��K �����X
�E6�W�X��%j_��%j_���`_
��M_��%1_�E6�W�Iu�T�l�����,��"�+y�lj��m0�'_z�'_z�)�{��|I���_���)yF;A�_��{s�_��%_��E6�W��Y�"�+y,{�R|���ѲgZz�_ۭ�R|���l���g�N��<�ە�vEu�T�Ku�$�S��M��K<����������g�,|�����Q�/���\�[�m�ғ/=��/���/����/�⿒w��^۞�� ���\�=G�ߋ���5�g��O�{oK�/��R�/��"g�+������K)>%n�x|J,����RɆ�J�����"�+yF7H��%D_��:_�E6�Wr���	,lV$�%���}	ї}	ї}	ѧ�"�Lag��/����/����/=�"�+y,;��|�ɗ�|J.���"A~J6=�ғO���`���%1_��%~���E6�Wb��O�ݐ�|I̗�|�����5!��+yF�б�>%7H��Ex�Wrn�Hj��{&���<�$�R�/�ܿ�KuϤs_D�%�eg"�}J���)y��3	�@~	�@~����X�7�.w�6�����r���s_��E���lVr�%D���/"޿?!!�"��+�qF��_�_��ғ/�ڧdR�/bٿ�d�I75�En��lJ�EH�Wr�6��R�/����/rӿ�7�@��W��~D��Sr~DI1�Jޛ�C��K��'�J�	�p!��+yF?ۄ�%�Q�4�K>%��_�E>�Wb���%_��%_�_�%�j7��/Y���/Y�"��+��4�K>%a���/�Ϳ���l>%[��|J.�Ƨ'_z�'_ğO�^H��Wr]�BBҿ�K�iN���鋐���l�d�O���:�J���K��W��
�u�B��:_��:_�%1_�E��Wb���:_��:_��E��W��䋬����l����/��"�+���|�ɗ�|�ɗ,|����{��!�_�[hg"}Jn��:�J�B��n{l>%���{����{I���{J^�=Gʽ�?�J�#�^$�%/���K�=%����%�^"�%�^"�EH�Wb��E��W�"�)yx;�n{J�h)��r/)��r/)��r/)��r/)��r/׿���Τ�^"�)y�n�HW�J�	��{����Rݥ	���{	���{	���{	���{J��]y�_�E�1�݋�����m����^���^R�%垒벉J�A�_�u�W�K�Ȇ�J�/7���%_$�%��h=��/���/��"�+�.=�ғ/��R�/R߿����J�A�_��C��Wr�UR߿��p��`_
��`_D��?�_��^�'�����G��WrnU�Ku>%a�ӓO�c٬o�J��M ��_�3�z��\}	ѧ��L���M_���M�����՗\}�՗\}iӷ�|�·,|�§�{A[��[�o߆�oY�|o���<#Ma�·,|J�?�����͖l�cK��e��'�z�mR���o�ڧ��YM�3�`�I�[u���ĺo�&�o����o���\*ߥMɥ���y�[����[�M}����s�
��`��oQ�6�}�ܷ�}�ܷ�}�ܷ�}���M}�j�m�6~�e�[F�e�Sb���-��2�-��2�-�ߦ�oe�6�}���[l?%o5�}k�f~��O���-���O�u�j�����m��6�}K�$��~+뷌~޾���X�-��2�-��2�-����ގix�6�}��>%�_�b�-��Ʋo����o���o3طf~J\�v/���Ʋo���o���oe�V�oe�V�oe�V�oe�T�<Rn��6�}���~޾Mjߒ�mR���o����o����o���oe�V�O�E؆����m��o�շ���t����������o׷JJ.���~��~+뷲~��Q�[3�5�S��6+����ưY��*lVag��O����O�;�/I�6~����~���%�[��%�[�����*�m\�V�o��V�o����o���o���<��I���S��F�ﷲ~�M}���m����o����9�/��V�O�Eج��[����[��M}������*�)yF�2͆������*�����o��V�o��p����|X4T~���������9n���[޿��ߊ���ߊ�����7�-�1���mf���o���o����os�$J�U[ڱ�	���]��i��p��$���~c�%���m��V�o��V�o��6�~J�ˍ�a�[�M��l��6�~J.�gQG�1������v.`�F�M���l�����Ҝئ�oG���������vT`;*�͙���O�˶9c�M�ߎls�9�ہ�)�q,�jKs�`;P�(������ˀ�)�T[Z����v^a��Ϳ���o����ه���v�a;���}��>lg�䝰�9!1%�gF�o�&�C�q��8�v�a;�t�:l�ﷳ�ه���v�a;���}��>l�S�d���va;P0%�_v9c���Nl��i�ہ��@�vz`P�(�l
�ہ�m��v�`;c�(�l
�����@�v�`J�B����I����v�`;v����N"l��c��m$�v�`���D�N"l'�����)�.wi����v^a;��N؆�o����1��l
��RmV�-�c�����v�`;v�;؎lc췓Sr]>xP�a��+l���
�y�)yF[��
�y�m@�6�~;հ��N5l��S۩�mf�v�a;°��N5L�E�Ҝ}��>lg��۩��T�v�a;հ���:l����m��6�~;!��؎Cl�!���l|�Cl�!�1��	���vBb;!����NHl'$�Sr��Zg���ه��Ô\���d���vBb�l���Ml�&��	���vBb;!��؎Cl�!���q����v�a;�t��gt����v�a;�0%a�ub��t�:l���۩���v�ac��W��+l��������va;v�(�NL�c����mf�6�~;���D��K��9��N؎L�u�@�6>'�ہ�)y��4#���H�m$�6��a؎0lG�)�۩���v^a;��۽�a�۰�)�TL�`��n�N�'l��3S�Xn��n���v�`;v�;����6'���I�m$�v� ��'°�0�>L�G��p�!L����d�p�aJ��6N5�Sa�}v�>����C8��>����C8��>������sK.���>���-yx�Q�TC8�N5�S�T���OK.�.�0�#�B8��+��
�B8���̒7����\�p�!�j�©�p�!�j�©�p^!;
�pz �G�Q�/Kݒ��Y9��s_P�%�c`���뇣�@(�C������p?��!����,�����?��ap~(�C��mYr]l����0q?�G�Q�pT �"U,�ې����@8=N��_f�%a�1�?(����p� �1g���ߒ���$B8����@A8P�IYr<?����A8v�|��\��4�±�p� |@8���3`��ݥ9v��c��A��������G\,y��B�±�p� ��3���l��.��p!�D'�I�p!�D_!�B |�@�
�p�!�j_!:�S�7g�옾���Ēg�c:��=p��t©�p�!�j�����C��p�!|�@����o[��B��p�!|�@8���ϒ��=:�0�s]�1}�@8�0%�k�1���!�q�p�!|�@8�:���C8��0�#6>��y�p^!�W��y�p^!�W_4�0�#Sr]n}A8�:L������c�C�o(�!�q�p�!�}_Z�C��Sr>�:�N5��1�A�p�!t�A�p�!t�v�>���� ��Sr���c/t�"|'B8Z�V���E8G�Q�s��C��p�!t�A�p�!�j_G:���TC8�N5�#�$B8�N"�cS��Yې/-_Z0%�B��p�!aG��L�u��r�!�j��y�)yx;�#�B8�� aJ�h[G�:�W_��&!|MB8�:�/Sg���ݒ9!NH��Sr�v&'$�	�pB"��!�q�p�!�}g�هp�!t������C�S�TC8�0%�㩃�TÔ�F�ri�t�!t��>L�u��o�'$·C���8D8�>����C8��>���K��7�����ܸ���)y�6Q_�N[���E8m��!�0��p�"��_�`�s�E8G�Q�s��D84�C��\'$�	�pbJ��}�/f'$�	�p�!|Ô\��B��NHL�E���&¡�ph"��'$�A�p�!�j_��r!�}g�ه)����j�&�	�p"�}_��C���8D8�C����C8�0%�hgr�!t��gt{��C���p"����C����C8���!��A�������L:��S�v&��:�SS��^��p�!a_�N5�S�C8��0��
����e�-ͩ�p�!�W���p8!�D'��7��j�±�p�`J��U�/'�I�p� ;_����@A�ʅp� (
��)���������FwVe�r� (
�p� (߯�_!;�±���
��A8c���Ig��p� �1g�w"�cS�mi�&!|B8�� !�W���p8!�1g·�o;�±�p�`J�	�S���;�w"��DG��p�!a'±��e
��Q�)y�n�|�A��)y�v��[~'�I�p!�D'�I��e
��)��
�pB�2��e
��)���C8�:���C8��0��
�B8��+���{���q�aJ��8N5��?�d���[�Sǩ���q������T����A���q�aJ.��w�}8�>L������q�)�z��;�Cg�SS�����ot��g���!����>'$���8M�&���q��{��}8M�!�ot8�C�!���q����q�����)���q�8�pa8�0��0%O=:��I8:��I8�.�;���ه��q�aJ�/g��D8�CL�uٙ�8�9�8!q��8NHL�;�7n�	�����6��qBbJ���8�q�8q�8�C߉p��8NH'$���q��8�q�8q|s�qB�8!q������g��yb=�_�8�p�W8�+��/@8N"_�p|�q^�8�pN8'���RmV�+���I8�+��oN8�0G�#����q�aJ�����TÔ<��k��r��8�p|M�F��#Ǘ)��/S����ʅ�+���A���q��������
ǩ��T�q^�8�p�W8�
�oN8�L�����Y�8vp;8�g��W8�L�E���p�_�+_�0%���q��8�p�W8�+_�p|1�q^����$�q��ʅ�+��
�y��+�#����q�aJ��^��q^aJ�����q^�8�p|1Ô<���w5����"��B����ۻ��	a8�0L�û%s^�8�p�W8�+���	�I��$�q�8�p�D8���;�vH��%E���7����jxO}2 )=A���*�]/�v5\�µ����*���b�+Nx7Ǯ�+a��kWÕ0\	Õ0\	��+\��'\%�U"\%µ���8�E�	��W�z�+N��+N��y.�
W�p�
ג�k�Ë<��O�p�}x���P!�"��b��M\�!����(���&��W4qE�*�y��/���g� �Zq5W�qm���C\�ƕi\Ƌ�x��U[\#���-���-���E���Nk%�L�Z+qe�Z�+Ӹ2���x�w�Q+Ӹ2�+��Ҋ+����k��M\��M\��M\�ĵV��(�h��!quWG�"�ꔓC�ȏ���*�+��
�+��r�yW}�TH\� �h�&�h�&�h�E�h��h�&�h�&�Mצ����:����:������qstWG�"��vb�ċ�l;W�q�WZq�WZquWGqu/�/����ZquWGquWGq-��Y\��U[\��U[\+*^��VT\+*�&�j2�&�j2� �ZQq5Wmq-���+���+��VT\M�`��;ጶ��E��d���d\[+^�7:D�!jE�s\��Un\��Un\��Un\�Ƌ<�sU�q-�x�G�Sr-Ÿ���������]���v�ZwqU W�~���Q}�s\��Un\�-����mq�W�q�W�q�v[\}��w\}ǵ��ZwqU ��+�+�6`\��Պ\a����!��+��︶V\�ǋ�F(%W��".HrU WrU W�q%W�q���k�ĕ|��g�
�ZQq����O\�U���QQrU צ����O\aȵ|�jE�V�jE�}W>r�#W>r��y.'�MW+r-����Z���Z���Z�+�+�kEŋ<�#M>r�#/�\�BE�U�\�ȋ<�SQ�"����\�.�81E&WQr-Ÿ"�+2�"�+2��]\�.����N���L���L���E^�S>r�#W>r�#��k����s9D����]\�-��/�>P�Z���ڀq�./�>P*]���jX^�e;+W�r�θ�+X���k��հ\���\��ǹ*k���+ky�G��Dm�6s\Y˵���Z^���S�J���+�/!k	YKhXB��Н��$D&�	aHCB*�P��
�E^S.���Hؓ�d��s1��P���$�1�B+Z�Њ�0$�!a�Fئ�Њ�V$�"a�F�G�?uC>򑐏�V$�"aOF�GB+Z��:#�#aOFؓ"���ț�H�ɋ<��k9��(a�F�NBw���Y<���ӋLBd"����$���H�GB>Z����^��ʂ��-	;7B>l�!2	�I�LBd򑐏�|$�"a�FhEB+�����}GX�6`��	H�@B�b��a)Ƌ<*?)CQ�"�3SX��b�%�(!E	)JHQB�R�P��!2	�I�LBd�d��$t'�;	�I�NBw��Н��$t'a�FHQB�l�!E��xT��!X	�JVB�����`%+�N	uJ���P��:%���J�S����#4,�a	ˋ<�O|J����5aGX�z��s#�/!~	�K�_b�xg�F�_B�����%�.�a	k8B�������%l��K(]B�J���#��k8^�_ =L�aBJ�P���%d-a�F�ZB��"�\U����ty�w¹*~	�:^�Q��z��Ä&�.�t	�K(]^�7�pj�G������E�q81U3a�GiBz��Ä��t	�K�ZB������5a�Fئ����`%,�uJ�SB�l��C8��O��а���a	KhX�а�`%+auFVB������a	K\��D&/�|�ӝ���E^��I�R����%�(!E	�I�NBw�"o��ʲ�Н��$t'�;	�I��R�y.�(!E	)JXꔐ��%t'a=H�v��%�	�@����*���$%/������$D&aH�LBdv���{�_8m	)JHQ�Ɛ�$�	KhXB����#�)!E	)JHQB���Н���E|��w��NBw�"��Y�N	uJX�����#4,�ay�Gu�SBw����e�;	�I�LBQ�u���EBQ�p��$%/��r�S���$%!	�:B>Z�Њ�0$T �	�4B*�P����E~��I����M#�a�F�;B�b�y痾#���}Gعvn�
�E��)��}G�;B�2��`#�a�F�9B��"/�)��x��r�Y�*�P���s	CB��0$�!!	aHCB*�P��
�E@�@B���|��#l�x����
$T �	�@B�"�����-�	�HhEB*��w��#����F�4B�j�y��_����#l�F�-��`��",�6B�j�P[��C0B��`����c��92��i�L#4��MFh2B�����#���FX�ʍPn�r#�aG�9B�ʍ�i�L#d��iEH+²�P[�菏����f�G�4B���`� #/��4MFh2BZ6sD�+S��P[��"����;B��P[��"�aG���`� #l�MƋ�k"��E��X�a�G0B��&#41�B�:BZ
�PH����1J!�u�e!�x��r~�(BG:��Q�B"�	�DX�
�PH�-!��D($B!
���#���D�!B�ڇ:��!,��:B�B�:��!�/���K�ڇ�>��!m�H[>R���s���\i�G�&Җ��Q���~��)�H�9�f��s#�)�HiEڹ�j�T[��"���HE�(RG��u��"EiGZÑ�p��"ui�FJ+RZ����s#u��Hŋ<3�����"�ypK�Dڦ�r��C���3�R!�
�TH�B"iG�!R��">~9��)�x���5.~��h"-�HE�ߑҊ�V����H�E�-Rm�j���#i�G������HMFj2R��"��Y����Y(�H�AȒv��r#)�H[>Rm�j��Y<��i�F
0R��Ҋ�V��"�)�Hiŋ�8���d�V�ȣ�Ҋ�V��?4��/�\Ҋ�V��"uiGJ+RZ�Ҋ�Q�h"��H�D*$R�r��C���J��B�:��i3G�!R�"o��_r��C��E�a��H�D*$R!�"O����Q��"u����OݔV��)�H�D*$R!�"��kS!��B"�)�x���1$i�Gj�⏔C�"�)�H9D�!�.���#��H�CjR��ڇ�>��s9j�/�������$�i�GZ��r��C�"-�H�DZ����M�B"�)�H�C�Җ�'�eiYGJR�ǻ��S	CJR��0�^!�
�WH+=^��;������hHjR��ڇ�'�O]�DZ�
��$E)�H�D�&R4�փ�� /⮪-�Ɛ`�%"��HF
0���d�&#5icH�4R��2��i�&#�IMƋ<�sU��V��L#�I�F�+�ʍTn�r#e)�H�F�4�^�y.�W�/�\>��@R���`��"-�HF�-Җ�`��)�H�E�-RG�:���#�)�HiEJ+RG�Vz��"i3G�!R�r���#��H�;����V����H�E��Vz��"�iG�(RG��w���E����H�EZ��j�T[��"u��x��壢���H�;R4���M�h"��HEZ֑:�y���"���H�?R����Q��"u��HE�(RG��|��i�GJ+RZ�Vz��"�)�HiE�(RG��u��"��H�:Rm�j�qsi�GZ�2���#��Hiŋ�FG�e��H�EZ��"?�B�s#���H;7�΍`��"�i�FZ��j�T[��)�x��RH�B"��H�Dړ��d�h"��H�DJR���"U�jHUC�RՐ���0���JR��0�?F���Q5��!��H�C
Rv[��)tx��p~���R�TH�"�)aH�� �P9�T/�|�*'��!UiF
���>�iFZw�"��H��"E)�H�DZd�Y�E)�HiEJ+RZ�Y��"�/���)�H�EZw�j�T[��)�H�D�!^�g9���H9ċ<��J&�H�D*$R!�
�TH�B"i�E�!R�"�ÖE)�H9DZ>�B��|"-�H�'���-�Dj^�7:���}H�Ë��N&9D�!R�B����!�(�>�TH�B")tH�C���0��!%iaD�RՐ��T5��!%i;D�Rv�����!mtH�AZ�<�� �oH�R��J�T"��)NHqB

RP�"?�G�A�Ү�T"�!�oHqBZߐz��+�ȣ��4> I�އT5��!U�jH�B�Ү��+�^!�jH[���0��C�oV��0���v�(J�PJ�����	%N(�J�Pz��+�8�E��e�C�^�x$+	C�Q���j(UC�J�P��+�^��
/�L��+�^�E~<�_eWCiJcP����4%((�@�J=P�y~͕]eWC��P�yTV�ʒ��0���,y(KJ�P��+�^��	�D(�^�e;��
�W(�J�P�q.UC�J�P�)�j(UC�JcP���T��3G=P�>�ț�������x�����%%(�F�R�z�E�h��ʒ����/�F;���x�z��p�-痄�$%a(#J�Pz�'�8���(�B�J�PℲ��
%;(Kʒ�R"����D���'���e�C��P���-%;(�AY�P��eC)��R"��4e�BiJcP���Ơ4%((�@�JP����.�te�B� JP"��&�t�(]@ٜP���9�teMB�^�7:�t�(@� JP"����Dx���%(@� JP"���D %(7�˚����D(@��_�����/��>l�vP��m�zYmPV�����cP"�yَ4]@�JP"��������F�,-x��谲��l((]@�JP��r���/7���d��~��_�ߗ���}�l_.ۿ�r��ܙ/w�_��;`\�/��˝�r�,-(����Ǡ܆/���m�r�܆/{�m�r��\}/���=�r��E^��Q���R{��^��=eiAYZP���eiA��^{��R{��^�
��ot��*P�
����6|�_n×��/���B����{��^������z��^������z�P.�����k�����	�l(w����r7��M/���"�h]D/��E����k�+|r��E�G_�_.������i�=�rϽ�s/��_�7:`�`/7�_�7���R{��^n����z�P��}/�\N9���=�rϽ�s/��˾�r���(W����r��\}/W����q.W�_Ĺ,(���rA�܆/���rA�܆/������{�ҹj�@Y4P�����e�@��^Ee�@�_v�{�e_@���r�r���(��˥�r���(+ʥ����4��=�rϽ�s�wf9@��^����e9@YP��� e@�F_�ѿ��v2�Y_n֗k��}�F_6���/W����rϽ�s/���W����/���=�rϽ�`/���u����z�����������{�/��e�R{��^����s/���=�r��\W/��˷��o�/w��E�r�E~�����r7��M/w����yT������y�u^n������e;�\W/��˾�r]�|{�O^.�����x�)^�^�\/�����ry�\/���w�����x�<^�8�\/�����j����/ߥ_���ȏ�9����������}�����y�O�"�4q���'/���w����7�i�y�b^����s9`|�~���r��E~�3��뗻��nz��^.�����"z�b^���/��������W○��������e��z���"�Hs��E�hߥ_�������r��|/�_n×���6|�_���E��$���m�r�E~���m�r�܆/���m�r���s/��˥�r���`/7�����C8�s���1����%��{��^��/W����r��\}/��_���\}oW����v��]jo��������R{���.��K��{����odb��/�N0���K��R{�^�vϽ]jo_���C�x�n����b���o�����������k���|�3����?_�F߾��}/�Y�nַk���Yخѷk��}�F߮ѷk��}�3��̷;�m@�Fߖ����f}[�.۷��m9@�ߖ����p�n���3����v%�]�oW�ە�qW�����h�]�oW�ۢ��h�-x7��v�-h@� Z�"�����.�u/�Nr�@�*����m_���ю���V�z��-h�Z=��V�z���x�w�Akڶ����e-;h���<��^c��^w�A�Zvв�����m�A[mЂ��z�E�^=�R���N9@�P�6�T�u�h]@[G�"����u�hKZ*Ж�z�--hAA[Z������-h������1h����_�B�A�Zv�"��HS"��C8���Dh�A[Gв����-;h�A��:�V"��;��R"��e-;h�A�=�J�V"�u/ⲕ-;h�AkZc����Ơ5/����h�-h%B+Z���E�Wh�Z��z��+�^�E��E��+��C���WhqB�چ�'�q��Z�Ж����
�WhKZ�������	�Dh%B�P�6�^��
�Wh
چ����m(x�Gu<�P�r����mCA�&Z���Em����F'���u��hE�(ZG������#h�Z���`� �m(x�GuF�4Z��2��i�L�em�A+7Z��ׁ��h�F�4Z��2����E~�Y��"���+�x������E�U�����W���������h1G�9Z��ʍVn��miA_�i���Ǡ�!/�\N_�Z>�򑖏��(iEIkEZ+Җ���i�HK>Z�і��-�h�ڢ�V��
�U �iH�@Z�*����E�ˑ&iaH�@ڶ��w��miA[ZВ�s�r��#h1G�9Z���������h}G�;Z��b�Vn��ot�����r�e��hMFk2چ��i�L�e-�h�F�4��`���h�Z��������x����B1G�v���� �%m�AK>Z��"����0�U �ik�N�֊�/�>�HkEZ+�Z�֊��i;^�e�\(2i�I�LZd��+��E&msBۜ�"���Ȥӹ��U+^��q�JQZ��"�娕����(-Ei)J[��R�����mth������5,mWC[���֝���Wh�Z���+�`�+-Xi�J�SZ������ۣ:�mah�JVZ���.��ж0���mahYK�Z��V��ҥ�.mC�_Z���y.'���0��i=L+]Z���Ĵ���jx��p����ښҴj�U3��i�̋<�SH�?��-�
�E�����i;1m�h5O�yZ��"�ѹ*�i�NKwZ��:��䡥;�>vJwڒ���(�E9/��}z�
��}hKZ���3�t��;��iQN���:�����;mDKwZ��ҝ��N�m�h�N�tZ���>����i�΋<��O��j��V�>��B�O�4��������hk%Z����V�5?��i�O�G�nwb��HeЋ��,��e@-jPk~Z��v[��>/�>c�yZ��Y����</���IT�Ӛ���5?-�i�O|Z��v[����x�w��B�NKwZ�Ӣ�yzg�N���h+*^�9>-�i�O|Z�������E��Y��i0F�3Y��g4?���,F4������g,���HwF��"��)7�Q�tg�;#���HwF���kȏg��}��+*F�3����g>#�Q΋�,���tF�3:���(g��QΈrF�3
�Q��gl���hkF"3��Ìf�0��=��aF�2�y�<ˍf�.�t��(]F�2J�Q���ed-#X��VF��"�����_����:e�)c��V�"�Ѱ��c��(]ƺ�yT��f�0��=��aF3�i����8��Q͌jf$2����(]F�2������#Ey�7�)�x�{�Gu�Yw1R���b�)c�ŋ<��O��"!X�-F�2����b,��ʋ�,��4,�G��w~iXF�2��ѝ��dD&�(E�(J�>����|d�E�(JFQ2��Q���d%�(y?��,'�0d����416M�����G�1�����	1ǈ9f;l�1ǈ9F�12��bl�� F�1��Q[��?������ŋ�xHI+FZ1Ҋ�V��b�����(F41�<�hb,y�Ĉ&F4�"��	����(FG1��M�b�CA1r����jM������(F41ڇ��a�c��hF�0B�:��a��� �*��C�U#t��F�0B�:��aT�jUè�*����`#(A�
FP�"���V����E~�cH06:�T`,yKF0n������c�È ^�!�9����.`t�����xg�`D #x��p2���"��7�Ǎ�q���������
b���� F�"/�ca�X1���bl����1R��
�T`��]���*����s9���#F*0F�z�EՇ-��X1�����1#Fc0���`������v�Q�U#(� Fc0����ca�(�Q"��s9D�	#N���Fv0�����`,��!�އ���`4�1��h^����`d#;��hFc�"�\�Vb#(A��<�sUP�"����#;���Fc0�Q��`d�1��hFP�"�����`����m1v[��`4�1��
ƺ����`4�1���F0�����k�
�T`�c�ŋ8��`#(A�X�1�b���E��Q[�Z�3���+�^a�	#NqF�0���+�^�E��:}�
SQqF�0ℱMc�
�W6F�0z��+�ȣ:�%#a��ˁ,a	�(F�0J�Q"��`��x���*�F�0�'�8a�	�D[>F�0�|�^a��qF�0�@���`dc=�(^��!���U"�a��D%�X52�'��"#Nx��p��F�0z��j�E�˧ZIF�0���aT�j�GF�0��0���rʉF�0J��Wd��Dx����g=���z��d��1��hFc0����`,��hF*0���d��]��F0�cJ��Q�z`����ƪ��.`tc�H�.���c,�]�� F0n����/�}��`,�]��F0�����#��HF*0փ�� /�>CFP0v��] #;x�������`d#;���Fv0�����`d�1KD^��U�(�W���|�2J�"��_�g���/�F~����"/��Y�����/
#�;1��C�>�}�w��Y�<��\�"��;W�������E����<����"��;���[�;��ȣ����/�?��ȣ�N�/���y�~���;��\�E~����/���y��g�/�\�s��<��}���"��;W��s���/�O�w�~�G���/��%�E��w�~����_Ĺ�su9W_Ĺh�"��8�/��@+�ȣ�>�~�Gu���"g4���F'9] _���E�hh�y2����F����y2�⋼l�/h��;�E5|�����E~�s��E~��c����U�����BT�����C8s����y�0�i|߸0�iN�"���E�U�4��ot(@��C����"ᜀ0|���v(й�E~�n؇/�l|�GuNЦ�E��7��y��7��y�	_�5����"?��w�yT��_���dE)�y}fBH|���ch�<��Q8�/�����"O�������?�?O���">�8� _�7�-�ȏw�0�ȏ�9������"����sr㋼����E�{g!��<����E�Y��x��L�d|��p�Q��E�� _�!��	��"���~��pB>��o���/���d|����S��yT'&V�EQ`�y�(0䋼l�V��x?R��E�i;�!_�!�!_�5�@^�,�||���E_�5B>��s9D)��"��x���<�S+�E~�#�E|���H�|⋼�>�aE��s9�����/�i �/��}����FG勼F��䋼�>��N��C8Ҡ(/��Q�"G%��㋸F��q�(�/���/����@n|��� s|����||��r�@>�ȣ�d��"���E~����E~����E^����E�hGU_�7:M�_�!�&������"摒>ȍ/�N��y'�&�C|�G�	��E�_�`�/�>l�9������<��d��/���U�'��sA>��sA>��sA>��s�O��Q|��r cE��C8�Q _��q�B>��;��M�/�/r�C��C8�i��"�@�|�7���V�<�c;ۈ�9�%_�Q���9���"���Ê|�7�GE��ys�� ��y�;_�wlC��;��Ɗ|��plcE^�@�|�<��>�E|#7Q�E�Q�E�E~�s�E~���E~�C��E�h|���x����E��s|������Q|��p<�;������_�7:��_��ϫ�J|���H�C��x�&㋼ �1�/rXA+��r~A+�ȿ&N&ŋ|����<�󋮆�G�E\6���F����"n��<��h�/��PG[|��p�0��[��C[|���m�"�⋼_N9h�y.���"��E���H��y.�#L�<����s!�_乜���/�>*R>�E�9����"��?P>�E�˧G�&��?G-
��F�!_�e;}i��"��@�i⋼�v�V��Ê|�y�?��_�Q���"n!��<���އ/����/��G��y.�#0�<�+�E�!
�"��ĤC�<�CQ�"'&|�<���X�9� _�e;Q _�7:��_�g9��_�]����"��<�?��}�"?�aE��y����d,M��d����v�/�=�Rn��C�Sw�4^���\�dK�����"/����Km�t/�̜��X:�E��yz�RH,��RH,��RH��;�S�RH,�Ģ
�<OiKG�tKG����"��ߵK4�DK4�D�އ/�y$[ڇ�}Xڇ�}Xڇ�}Xڇ�}XF|�7��K!���v�/�\r�%�Xڇ�}Xڇ%tXB�%tX�E;�q��%aX��WXz���^��PհT�v�/򲝅z��WXz�%NX�E��y�N9���C8��K谨ox�Sn����o�"�ё��_�'�E1�y�VB�E}�y��_
�E}Ë�Lr�E}�y���c��ai��ai���+'�Xr�%�Xr�%�Xr�7_�FǐB�E�1D�Ëڇ�}x��Ö�aI�^a��^a��^aQ��E^�ӄ��/����䜐0,�ȏwtP��E~�OC���jx�7�#tXB�%tX���jX���jX���jX���jx�GuX�4�E���t)$�Bb)$}_ĹD/�\��E�ŋ|��V,iŋ<��OZ�tKG�tK���K���K�h��"�hU���$aX�E����>3I���E��g&�¢���,��$K��?��?Z�~��^a��8a�Z�"��q2i}_乜9�E��q.
#���ⲯ?��K*���v�/�}���C8��>R��q�~I�T`Q+�E��!(XꁥX�J|�Gu�\g��`i��`i��`iE_�Q}��N&%�R",�.��s��:Ү#�:��
K���
/�\�4	Ò0,	��+,0��k���R�/�|4`|���c��du}�RH,9ĒC��C($�Bb)$�_乜�:���X�b|����J4�DK4�"��!*�X��%�Xᨥ'㋼QJ1��otbRw�E^�SN���"�/��*��M,��
��_�g9�DK!�K��K���K����n�/�N��]ڇ�}Xڇ�}Xڇ�}XB�%tXB�%aX�V|��0,	�'���',q�'��C8��
K���
K���
�֊/�\�B	Ò0,q�R",**��ot���^a��^a�E_�Q}��+,���+���P��(��"�щ)NX��%;X���1X��1XTT��Г,**�ȣ�#���/�\�Uq<�sU���	K����x����x�,��R,����⋸ �'��o�h��"?�)G����N9A��0�<�#�/��4���
,z^��,z�ȏ��M*��K�tK�t���/���UP�KP�"��H���s9����/��L��1X��E1�y0����-����EBP�KP��K=��K��1�>�I�T`I�T`� ����/��!�j���_n�/���������.�r��˿(S�"o�#������rq���\����e;���y����J�r%��ܿ_�c�_�!�_n�/��]_�i.�/��]_�p����ܿ_��/����/���r��tK�E�{�����F�/���s��޿��_.�qX���\�_.�/�����R�����_n�/���[�������r�~�Y�\�_��/��k��/��_.�/���_��Q�>���[�˕�E1�yTg�8�YH}�y|��/��������/��B���s9�j��?��-t�J�T�Eչ�X�yT窠`
��`���[=��ClA��
�E���v�-;ز�-;x�GeFo%<*c{[�-��z�y����-a�FlUöb���a��U[հ�}�z��W��m}�'��odlo���+l���+l��9���VA�ȣ2���a���[��mt��m}Ë�F��V5l	�'lq�'lq�'lq¶�a������-N�ℭDض0lq�'lq¶�a�°%/�N�^���'�yz'��ak��[��[���[���o�ڇ�}�6:l9Ķ�a+$�B�E�˹�}؋'�}�ڇ�}�B�-tؖ<lK�b[��/�\Q� �hb�&�hb/���a[�Uے��jؖ<lUÖ0lK^�5���"�b�!�b�!�v~�!��a��a����[谭��ڇ�}�Fl9ċ�9N&;$��b��E[4�E�w��/'��-���-���-��j�-��Ҋ-���Jlk%� c�-^��{{[+�5[���[m��/�����-���Jl�`l�`l�V[l��V[l�ŖVl��M��C�(��b�(��b�G��[Z��[G����ҊyT��q�
0^�Q�2���ضVl[+�Lc�4�[����>���x�w�Qk��wl}��wl}�Vnl�Ƌ�x6[>��/���Q��*�-���������mEŖ|l�Ƕ�b�@^�-tF�Z��"�"�mkŋ<�Yd��غ�m���l[+���֊-E�R�m�Ŷ�bV�e[w���xO>���۲��a��m��ְl�ְl�ְl�-�`�E�	'��ekX��ekX��e[��5,[���)[���)[���([���(/�~���;ٺ��;ٺ��;�"�-2��dl��֝l���l���l�ɶ'c�N�=۞���ヮ�ekX��/��ZYˋ<��کty���AW����-~y?�8�f�a�f�_��e�_v8��/[鲕.[ֲm�6�l��V�l�A��e�Z�-[ò5,[ò-���/|˶�ckX��ekXv8e-[ֲe-[ֲ5,��m�Ƕ��E~��Q鲕.[鲭�◭tٶ|l��V�lY˖�l[>��e�Z��e�Z��e�Z��[ֲe-۲�mY�V�l�˶�c+]��[鲭��◭t�J��a��y�1e-[ֲe-[ֲ5,�΍m�Ɩ�l���ȏ���:e�S�:e�S�eKQ�e[��m�غ�-2y���5:���؂�m�V�lu�V�lu�V�l�.��d�N��d�N�[w�E&[d�E&��mƖ����N����؂�muƋ<��Ϟ�mO�V�l�˖�lY�ְl{2��ekX��ekX�=�i��-kٲ�mu�ְl�3����-~�Vgl=���l�3^�Q��ll!��l6��fkk^�Q�r�-��6sl�V�l�V�l�͖�l�͖�l�͖�l�̶�c[��"?��,��f[��6[[�"?޹jǖ�l���l!��l�:��fkk��f[ֱ�6��mǖ��vb*p�g+p�g+p�g[ֱ-��:���y���7�Ng�t�e۲����6s��s91u:[��8ۂ�m��V�l�V�l΋<���h�ƶ`cKw�tgKw�tg۹����j�m���l5ϖ�l�����C8ۇS5�V�l�9��g�y��[�>[ͳ�<[ͳE9{���xg�(g�r�(g�r�8u:�΍y�tg�Sn|ƴ�ck~��g|��[��u:[��m�ضil5ϖ�l�3��[೭�x�7��;���l��V�l5�V�l5�V�l5�V�l5ϋ�FG�Ng�r�5[��u:[��8[��8[��8[n��6[n��6[n��5[[��5[[��4[HsT3��c��Q���Q����Yˑ�Y˱s�(]����Z�����qd-/��s<6s�Ѱ�̯#X9�p˱����q�.���t9�p����Ѱ���6�:�E^6��hX���΍#k9���a9��a9��a9�p˱s��Z���V�`�V�mG�rl�8��qˋ8����Z���S�:�L���,G����G^ğ�GdrD&g9�%GQr%G>r�#G>rl�8�i�4�mG>rl�8���(9�#9Z��9#9#y�����Y<l�ȋ<��j��"��H���X��"�ꔳ����q��8◣t9�w�ˋ<��o9�$2/�\�G܄4GHsT3G5sT3/�\����9��c���{E���hk���E��B�̑��̑����>*Jd�U#Ǫ�#�9B�#�9�#�9�#�9�#�9�y.g�%G5�"����hm���m�Ҽ�?4Ƕ���m���hk�}'Gns�;y����.�9��#�y��бm��Q��Q��+P�(�(p���wrD9Ǿ�c�����͑�m��;J�j�f���_��$G��"�ѹ��9z�#~9�cG�Q���Q�������Q��ˋ�N��S�}'G5s�/G�r�.G�r�.G�r�;y���,��=����Q���Q��ˋ<��O�r�/��9z�y.��X�r�0��c�ʑ��̋�87G5sT3Ƕ�#~9J��t9J�c����˱���a���_���_�.����y�ɛ���=���=̱��_�.G�r�.G�r4,G�r4,ǆ�c�ʋ<�C�:�N9���N9V�)ʋ<�SN�r%G>r�#G>r�#Ǣ�#9�y���)M>r�N9�#y�%�͑��ȑ��ȑ��ȱ(�؊r�!/��L�9cmɱ��@���H>����drl29#y��ъa��aȋ�F�0��wr,79*�y��WE+P�
�H>����wrT Ǿ��9��}��w�L���H>���H>����drT �ڒ��8����86��ǋ8�
��wr�!/�jE�V�hE�0�X�r�@9�#9�#9�yW�����(9��ȣ�SWdrD&��cQ�ѝ�R���L���L�(/��Z)�ѝ�ȣ:}�)�
��N9ꔣN9ꔣN9�c�ʱN�hX���hX�`�V�u*/��hYˑ�Yˑ�Yˑ��T���(]���(]���hX���hX���V��E�^w�?>��N9ꔣNy�h������R���L���(J���(J�V�@�
�H>���H>���H>���H>���H>���ذr$G�q�/�\N9�Ǳa�E����X�r$ǆ��9*��9����s9��a%9Z�c[�ъ�Y^�!�L"�#29���(9���(9���(9�������QQ+r�"G+r�"G+r�"G+�"o�CԚ�#29���(9���(9���ȱ����r%�2��>P�N��0�~�#E9��uʋ<���#X9��#X9ꔣ(9���(9��ce��E�Q�Eɱ�(J���(J���(J�|��G��0GQ�"���+c^�|.l�����"s��9ꔣN9���ʱX�hX�]3G�r4,G�r+/�\�m�g���(]���Eջ�V��˱��_��5�ޚcI���������l���(]^�!���=���=���m���a���a��_���Eձm�ͱ��i���f�j�Hd�U6�ޚy'|BV��̱��f�j�f�j�f�%5/��h�g�j�f��3/���W5s���B�+�����׮�k�̵k��m��2W�s8Wn�"��v�\Q���\m͵��m�e0W[s퇹r�+��r�+��V�\m���\�a��0WHs�4WHs�//����+~��+~���+k���\Y˕��ȿ�L�k[�U�\Y˵a�jX���jX���E\�`�
V�+׆��a�֩\�T�u*W�r�)W�r�)׾�yz'�:�S�}'W�r+W�r�;��k�հ\˵��Z���jX��(W�re-�V��t�J�ysxf�J��,��s9�d-W��u_y~�^��U�\�˕�\Y˕�\˵��Z�re-׶�+X�ꔫN�ꔫ;����;�V�\���\�ȕ�|�BF�UE�U�\Eɵ��Z����yz��t'WQr%WQr�#W>r�a����(������F�q8��!ߋa�<���V��5�F�g�L�ڊreW�qeW�q�WmqmE���\M��d\��U[\��U[\�ŵ�
0� �
0���-�E)W�q�@����ɸV�\�ƕi\�ƕi\�Ƶ��Znr-7�������+��ܔ�����r�+��������w\}�Un\��Un\�ƕi\�ƕi\�M��&������M�q%W�q%W�q%W�qe׎��ܸʍ�ܸʍ�ܸʍ�ܸʍ�ܸʍ�3��>�)7�M&W�q�W�q�;���+�b�+�b�+�V�\+P�����#�e�U�\�U�\�U�\����m�|T�\}��w\�N����;���9��&�r�+����+��GuFۊr�"��yTg��(W>r�"W+r�"ע�kQ�U�\E�U�\[Q���L�(WwrmE�R�km��\kK���L���L��%WdrE&WdrE&WdrE&�ڒ+2�v�\���\�ɋ8����Qru'Wwr�-y��&�+X���+X���k���\�ʵ���drm2���k�ɕ�\Y�հ\��\�ʋ�xG�`�
V�:�JQ�%׎��N�֖\�����s9�,7���\�հ\�հ\˵���Z��&W�r�;���\�˕�\Y˕�\Y�հ\�L�M&W�r-7�◫t���+X���+X�ꔫNyw�r��a��+X���+X���+X�ꔫN�ꔫN�V�\�ʋ<�S�r�_��kwʕ�\˵N�Z�r�.W�r�.W�r�.W�r�.W�r5,/�l!^�հ\��\)ʕ�\�R����N���E^�?��)Ww�`�F'���jE�V�ڊr�#W>r�#W>r�#�
��(���\�ɋ�F�N��JQ����N���L^�����~�SN��?>˻�ҝ\��՝����r�k�ɵ��jX���E�a%k���+k���+k���+k��kmɕ�\Y˵���Z���jX���E�����|U�\+P����wr�0Ws�0Ws�0Ws�/W�r�/W�r�.W��"��!�t�J��t���+k���+k���+k���+k��\��U�\��U�\Y˕�\Y˕�\�հ\�հ\�����?��(W�re-W�re-W�re-W�re-�ҕ+k���+k���+k�V�\��U�\{X���Z�r-]�z��t�J�kw�U���otԶ�z������\�̕�\�S���E~�CT�r-J���+k��+X���+X���+2�v�\��՝\�S��JQ����N����N����N���*J���*J^���{'��"���Z���v�\�S���*J���Z�rE&WQr�#�:��(����(����(��k��U�\E�U�\E�U�\Eɵt厳PQr%��+2�"�k�ʕ�\��Պ\��Պ\�S��)WrU W����;%�Ny��B��0$lX	�HC^�72���w��#�a�Jذ�"/�)�"o4��E��Y���#$a�J�@B�v��E)�	ȋ�F����*�!a�ʋ��L��t%D&!2�L��t%%/�������+����`%�a	KhXB��а��%4,a[KX��"�x|�P���%�a	�K(]B�V���%�/!~	�K�_B�ּ�&�ty��r�.�e0��	mM��r�yTG�'8��	N(p^�Q�	r��ۼ�s9�E9!�	QN�m^�7:}�4!�	�LXB�҄�&l�	[dBnښ�ք�&�4��	�aBHB�҄�0��	mMhk�~��&�	N(p�ʘ�('D9a?̋8�N',�	�NX:��&,�	5O�yB�j�P�t'�;��	QNX�"�?���'��	�ϋ<��W�v��('D9a�KX�:���%,p	�Y����%�<a5KX������m-!
P��2���%�a	P��j�P�+!�y���a��	N(pB�
�q����8��;��	Q΋<�cH���P��'8q�9
��a%D9a�JX�
��a�E~���-]	�N�tB�:����E�G��'�;a�JHwB��"�C�t�E�/��yB�ҝ��t�E��Yx|���'�<!�	�N�rB����('D9!�	KWB�:��('D9/�\�Z{XB�:���(�EB��"�Q�V��('8��	N��
�P���W��,!�	{XBnr��ք�&�5��	�L�fB5���ȄD&$2a�JHdB"�����E~��J�J�P����E~����H&k	YK�ZB����N%�.q�y*~	�K�_B�����%�/!~	KWB6��&�.�t	�K(]B��"�	��a	ˋ�F���_��D�(~	;]B��"�唳�%�0a�KHd^�|���%�5aL�mB[���ȣ:m~	mMhkB[ښ҄�&�y���!P[��P̈́j&T3��	=L��z��Ä&�.!k	YK��J���%,p	=L�aBz���%�0aKVB�R����%�(!E	�SB���Н��$t'a�JHQ^��qʩSB�R����%t'�;	VB�R��a�E��`%�S	uJX�֩��%4,a�JX���а�`%�N	�JX����%,J	+PB�������C���t	YK�ZB�������%d-!k	�SB��а��)!k	YKX���y.��_^��◰t%�/aK(]B�����%4,!X	{XB�����`%+!X	�J�S�:�Н�u*!E	�I�LBd6����=ky��LBQ��y���$D&!2	�I�L^�Q��������+�N	)J�N^��ѝ��$%�(	Eɋ�F�ɋ<�SN�v���$D&�(	�RB+��D;��#a�ICB*�P��
$T �	H�@B*�P��
$T �	H�w*��|D;�@	+PB*�P��
$$!��GH>B�V��(aJCB��$�!!	aHC¾�Њ�ț�od�H�G¾���$�;	�I�LBQ�����M&�(	EI(JBQ��P��M&1>�NBw��y.��%�(1����$,7	�MB����`%+!X	uJ�SB�V��`%�)�N	uJ�SB����:%�)�N	uJ�SB�R���$�)�N	uJHQB�R�y.��8�mE	[QB�J��(�E�ާZ=L�a¢��(%,J	�RB5��y.�}�fR5���Tͤ+)�I!M�fR5���yT�[!mXIVR[�֩��&mXIN�mRn�r���stڝ�����Y�Uftjk҆��֤�&�5i�J�mRn�"��M�M�m�ҕ�ۤ��E�e��7U3��I�LZ͒B�Ҥ�&�4)�I!M*]R�J�����k�y5-pI�K�_R��"/��ڴ&%2)�I�`^��4)�I!M�fr9�$2��I=L�a^�7:�$2)�I�LJdR"�6Ҥj&U3��I�L�fR5���TͤD&%2i�L�aR�z��ä&�/i#M�H����&U3iIMZR�ښ�֤��E�gߔۤ�&�5��ImM�[�ښ�֤�&m�ImMjkR[�ښҤ��E��I.�I�K�_R��">^�J�T���%�.)kIYK�ZR֒��T��:%m�IuJJQR��"����NI�g^�!�rvͼ�C��h�L�Z^�7:�SN���ϼ�kt2�H�������%5,i�L�N����~&�)�NIuJ�S�ޚT��%�I�fR���Ϥ�3/��&���`%+)XI�eR��ˤ`%+)XI�J
VR���ä`%+)XI�JZ�VƤ:%��I�J
VR�������E��G2[dR��R��X&�)i�L
VR��������$u'�;I�aRw���y'|����%�(i�L�SR��ˤ�2�aIKJQR��R�yǣ:%�)�NIuJ�S�~�ԝ��$�I)J���ä�$u'�;I�`R��R����%�IuJ�SR��VƤ`%+/��� �N_�e���'~I�K�5�����2i�LJdR"���2&�.�ty�����%m~y���\�äe0)�I�aR5�"�����u�Z�ښy.���2i�LJdR"���ȤD&%2)�I=L�aR��T���/�tI�_��T���%mkI�Z^�9��0�tI�K�ZR֒���%5,i�K
VR��v��`%�))EI)J�NRw�ּ��$�yy���_ܤ(iLZ�����`%m~I�J�S��y.�P�\(XI�JZ���T��:%-pI�J�SҶ���%+)XIuJ��I��R���=,i�Jڰ�6��:%-]IKWR��6���s9��))EI[QR���T��:%�()EI�I�LRd�"���$u'/�}���$%/��L"��%�#)I�HZ��Z�T��ȣ���&��|�M&�IH�;Ȓ֖���E~��D��"o�?U �yG��0$�;I�HjER���ȏw�H>R򑒏���E^���
�y.�V$�"iQJ�GR>�����$-JI�I�LҢ��%u'�;I�I�NRw���ԝ��$-JI)JZ����E)�aIKjXR������`%+iJ�S�
���`%�)�Ny�����$u'iJ�NRw�����$E&)2I�IZn����%u'�;I�I�NRw����V$my'%i�H*JRQ����#)2I�GRw������$E&/�N8�%)I�H
C�ƐԊ��C8��#i�H�G�^�yǐ|$�"�I�H
CR����#�/��>�I>R򑒏�w�� ��H�F*7�Ɛ�b��1$���H�F�4R����`� �E�a%�HF
0�S��p2�����d� #��H�E�(R!�~cxA�9D�!Ҳ��C�"��}H�C
R萪��0�^!�
)NHqB�R��℔�� ��HAA�̑����f���Ơ4�1(AA	
�f������e3G	
JPP�w���E��aU�w�ȏg2�����(�AY�Q�w��%N(qB�J�PJ�R"��%Nx��`�����D(�A�ʖ�R"��,�(�?J�Pz����)UCYRB��0���$%a(	C��Q�|�-e�G��Qڇ�>��sy'���j(%B)JvP����Ơ,�(�AY�Q�u��4%(�@� ʍ�r���/�-�-����E^�3���rq�\�/��"�rK�E^�c���rq�\�/�����r��l�(���e�rپ,�(���e�y�W����rپ\�/�,���r��,�(W��n�r%��(�-�"�r��\�/[+�]����E�ˍ�q.������Ȣ��/7�ˍ�r�l�x7GP���(]@YdQR��Ȣ��(]@�ZQ����E%(�@IJ*P����.�l�(0�����/��U�A	
J=P6`�eFـQJ���Ơ4�1x��Oݲ��E~��QvP������E^�Oiۉ)N(qB٦QJ���=�D��;N��H��Ơ,�(�@�J=�"O�㝠�,�(K1JvP�����d%;(�AٓQ�d�8��	%N(�3���+�^��
%N(�AٓQ6`���e�E)J��"����D(%B)J�PJ�R"����D(%B)�6��M�l�(�B�J�P��ۢ4%((AA	
�n��ۢ�x��p

JPP���T�D %(7��������5��/�,���r%�\�/W�˕��'�qq���_.�eEE��_��E�.��_.���~��_n���/��9v[�+��J���F��=eOFY�Qn�������_�����eF��_n������_�]���z�mQ���E/��(@� ʍ�r�l�(7��n���D %(@� �n��ۢt%([+JP����%(�@I�֊�
�T��%(�@IJ*PR��
���(�@YwQ���e�EiJc�"�����=eOF�*�����+�8��	e�F�*����s�E���k�FIʂ�R5���T�j(�4J�P�:���Te3G	J�P6s�5%t(k8J�P��0��j({2*���R5���T�j(�3J�PB��M��e�F�!JQr��>�ȣ:W��(�D)$ʂ�M��/�㝅:��Q�%�(6JZ�"��O]�EY�Q�`�ڢl�(�E�-JmQj��Q���t��x�V�����(�EI+�΍�s�E��j�R[�ڢ���(k8J�Q�`���E�G� �EէZ�E�-JZQVz�h���(�D)$J!Q
�RH�B���(9D�!^�!�ڇ*�U���RH�B���(�DY�Q��M��%�(�;JGQ:��Q����x��rԪ-Jm�"�QmQj�R[�ڢl�(�E�(ʲ��Q��k���,�(Ƌ�Fǣ&�E��h�G)7J�Q2�yTg� ����(�EY�Q�`��e3G	0JmQҊ����eYG�(�f��V����G�ot�	0J�Q6s�ڢ��(;7J�Q��y�i�u�L�4��(k8J��"�8|.�s�4e�Fi2J�Q�i�=%�({2J�Q��`� �,�(MƋ<�3G��"�󗴢�/�}�Ī-JmQj�yz�l�([+J�QVT�&�4��(MƋ�Cs2i2��i��;�s�}%�(�'J�QF����(�FYQ�C�L���(�F�4Z����䡥m}C���j�M�B�E~<?�b��Q��-�hE�(ZG�:�y.}ZG�:��ѡu��x�����mth�ZG�:��Q���E�	�c����h�E�(ZG�:��Q���E��h{Z�r��C����h�D+$Z��ڇ���b��>���-yh������E-�h�D�&Z4�v5���umWË�xG�-mC���:��_��m�B�-�N�� �E��1$�hiE�(ZG�:��Q��m'B�-Zm�Ҋ�V����Dh�E�-ZZ�V�ڢum�AK+ZZ�Ҋ�V���m;h�EK+ZZ�
�VH�=-�h�ċ�F��h�-@h�D�!Z� �B��Dx7G4�
�VH���/����r��C�С�mMBkښ��C���ms�9�~l�D�!^��ۧ4�^�!���(�h�D�&Z4Ѣ�M��max��rb���:�M�h�E��3�h�mC�&Z4�"�����V���u��h�ZG�:��Q��s�Obm�CK+�އV[�ڢ���hZ������5��h� Z��VA����h�F�4Z��VA�r�e-�h�F0Z���V[�ڢ�-�hiE��Ҋ�V����}h�E�-^�!|�<QE���Ҋ�Q���E^�SN�Ъ�V5�-�jhUC����+���r	�2�:����Ih�C�2�:�С�-th�Cۜ�ڇ�&��m�x����6h{���C�=��h9ċ�FG�B�E�ѡ�h�ċ�F�B���hZ4Ѣ�M�h��1x���/�듕��-�h�C^�]u�Z����0����
mi���lKZ��"a�A�^�7:�T�jh�Z��V���U/��!	Ë�F�s�ɤWh�B[m��y,JZ��z����e-(hAA
ZP�����E -��qō�v���o7��]�v���x�7�1���P�n����m�@��߮���/����s��߮�+���}�������}���E�����M�s�cA[4�n�[�����FG�[��~���n�[�����>����n�[��J~����+��J~��>n�=�~���n�[����������~���.��;�r%�]�o{����Ǡ]�o���5����ݬo7����v��ݙow��:�vg�ݙow��҂vg�--h���5�y.G����f}�F߮ѷ;��|��6����6|�=�.ȷ�m�@�=Юѷk��}�F�"�S�5�v��]�o+^�7:�\�o���vA�E�{�;���|�3��̷;���|�3�"��,t��]}o[�m���NL�_����tg�ݙ����5�v��]�粴�ݬoK�5�v��]�o��_��;1݆oW�������]}o
��vϽ�s����r��]j�v2Y4Ю����m�@��v����6|[4���C����v�݆o��ۢ����^�c�m�v�]}oW�������]}oW�������E���|�ߖ��|� �.ȷ��Fx��1h���5�vg�E���}�F߮ѷk�m�A�Y��̿�r~�3��̷�mi���F���/�\>�����vپ]�o���e�v������v��v�.ۿ�;��s��ݬo���5����]�o����ڠ]��q~�3� ��/���9��;�ci�XZ0��;�c���3?.ȏ����<=�>�R���>�����oVc9���>K�c���>��K��R���>.��K��R���>��� �R���>.��K�c������C0:�=�y�ɸ�>��?����q�}\}��r�qA~\����y.���qA~�s����q�}l�������[�����>}����Fj�=�q�}l[�m�y��uc��F?�яk�/�< �����l?.ۏ�����F?�̏;������_�B
�5�y'xf���e���`�6W�Ǖ�q%\�W�Ǖ�q%\�?;<�C�-�qK,@�]�qq\�����qK��{��qq\����-���`\��Ƕ�qq\���r o�]����q���w��]�qK��W�Ǖ�q%�1{�����`\�{��q%\�W����q�~�#���e���`\����҂q�~ܬ��e�q�~l(��_�e�@iC��3?��k�����3?�̏;����XG0.ȏ��/�.ȏ����8�q��F?�я;��6�XZ0.��q~� ?.ȏ�c���3?�̏���� ?.ȏ=��� ?6��c��3?�̏;�����P0�яk�/�o��ϝ���`\�K�8�,-K�5����E~���:���`�#�ƕ�q�~ܿ�����9N9��_��;����-�qK\���-���`\����-�qK�SΕ�q%\�W�_�!���Yhi���FG�[�ci�\�������Xm0���/��;�l;��Ƕ�q���w��]�q���w�Ǖ�q%\�W�Ǖ���`,-�밺�����c���<�#͍��q.o��k-@F0����`D c��� Ɔ�q�\�Kƍ�q�\�{�҂q�\���������E�U7����q�\�����q�l(�����q�\���r��c0"���?ܤc���c0���s9�4c��Xm0J�Q"��`�1%��c0��^a�1	�H^�]�QQ�0��m�}��hF�0B��0�c����0�u�j�^�!�c�XG0
�QH�b�c��!F1���a�
�W[F�0���E^�C4�����B���F��"��)'N[F�0z��/`�
�W%��Fv0�����o�N8���D[F�0�'�8alx���ɔ>��0�L:���}��X!0ڇ�>��aʑ&�9��!F1r��h`,���!F1r�:��a$#a� F�0���GEU��0B��	`��}�^��}��C�� #�9�h^�!�r��B`��jUË�,'�� �}x���5:��}�èF�0��Q5���E�ˉi9�X0���aT�jq�F��`4�1��?��i�|��(Fv0��������W��������7�a|	����Μv��F�0�'�8a�	#NqF�0�����W�<��J�0���	#Nq�>�IF�0�'�8a�	#Nx���)ͷ��8a�	�D%�Q����jFP�"n��`|{��Fv0����o���hFc�"o�OV�dǐ�`d#(A�
F=�"O�s��`����GP0��y'�L���/�_�?J�Q"�a4/�\�4_�?J���#Nx��ί��w���C��_��0���UèF�0��y.�}�}�?��
�/�F�(�Ҩ����)틖����_�~'�y'~'�����w_�e�N�/���C���/�G�y�ߟ�/��_�7�>~���;D_��c���߹�E�w�~���;D��s��/�\�C�<���/���E��<���"/�wb~�B�C�<���"��;W�ț����E��w���w�~���;1��o���_�!~'f������F
��?0������_����s���Y��"7��kt��9����}z�"��x�w������/�NL��yT'&��<��o�/�� �/��>L�y������"��Y��"����d��Y��"?�Y���?��;�,D[|�h�B��yz�#�	/r<R��E����"o���JL�q�0_�Qa_Ĺ0_�Q1/���E��^���NL����>*B+���;�_�!��h�/�| |��p<�-��?Z�( �E>c0��;�\�d|��r��4^�\En|��˹���"���s��<����/�?�ȣ:��W�"��@�L��F�*
���ߟ�/r��ߟ�_乜�(�/��U���C`E�����"�y�?�)S�"�\�Lዸ_�]D�yz�}%_�Q�X�/���X�/���+|���@Ɗ|��ޟ�(�/��(�/����K��ys��(�9W�!_��;jia�"o��>�"�(-_乜���/�\���\=�U��y.G-���F�*�<�sd�E�q��v���;�"�;�"��_�!���*�/򳜅4:��_��/�}8�|��pR�"�#��<�����/�\NL�ɋ�� �/�Q(�ys���;�"?��2�"o�S�:�@&_�]���v�9�(_�e;q'_�7��Q�E~�S��/�iX�/�����cE�����E�	Q�"��"_����|��*�/�\N&`����pX!J��;���|���)>�E|�ڎ!`�y�0�<��rX�/�+��yz�7��yz��G������"��xĊ|��r<bE^��C�|���!�E|�w��H��������|�w�(�"o����/�N_���q.���8��8��Ed����N_
6��;A�Ƌ|z��|��rF�3��E���}(}z���<�c��/�\>=�Z�ȿ&Nr�:�ȣ:ɩ��"��F�|���@��㋼l�*_�7:j�._�e;W�gLX�y'&���F�*��E������/�\�U��y�*����p��Z��o�|���E\6e/r<R��E~���EI��yT�(e_乜��u|�����"�(��<�C��E��Y�N�"O���s�<�#��/��>cV�Ȼ��m�y.`勼9���|�������/�\�Bˋ|�/�|�/�>�:�ț�%��<���~�"o����/�\4s|��|���|����l�c;i�x�O���/�|Tz|������|��r��m�ȣ�\�>��n�E���/�ù
�y�sn�E~��[�E~�[�E^��ʁ4_�-�)���/��/���!�9�ȏw�P��E�΍/����"�c����?��˦s��F���i�t�"�ч-���	��E~��d��/��q�I	~�"�����"/��A��y'��	�y�Oi��/����"�E�/��<�ӄ�/�\>�Ad^�dB�|�����E+��y�>l�_��C8�._�5���N��ߏ_��^���,)ʒ�,)ʋ<#m�S�:e�S�:e��E����1���eiX���E��[�E���Y�X\�E���'�x\�x�YR�%EYR�%2Y"�yz�Ւ�,)�ҝ,�ɢ���F�Т�㋼ ��k�G��c�9^�52'_��3M�rc-�r�E|��c�9�_���w,j8��s9'$K��K߱�K߱K��K��K��K�����"/��E��y.���rcѦ�E�i"�X2�%�X2�%�X2�E��y�N���d,z2^�ϭ%�X2�%�X2�%�X2�%�X2���X����X�EƋ�r����X����X��y�|��Q,�.���M�a�5�(^�e�m�E�)�}�>�.��C��C���-�X�%�X�%�X�%�X�]|�G���cqi2� c	0��bQw�E�	~.�`,�`,�`,J1��C�o�&�hb)$=_�pbғ�E^��Q4����?!���QG�(��"��ĔV,i��Q,:7��s9EK!�K���KհTKհTKհTKհ���"�ғ�E���|B�yg��aQ��E�/g!�_�Q���Y��X�i|�G�QQ!�K!��i�otg�b�!��a	��a	^��]K谄��/�:�$K°$/�N�H��y.G��aIm_��c��x'aX�%ax��0,�4��s�/rbҦ�E~���9�/��B��R5,U�R5,UË�F���a�=_�7:�$K°$K°$/�}�S5����񎂍�oi�'>
6��s�x'aX�%aX�E��y'���i|�G��O���/�>�]G=_���ঐx����b�DK4�D�΍/����}Xڇ�}XTg|>ޅ#M4�DK4�DK!�"�#M!�K!����/��8�K!�K!�K!��KհTKհTKհT�R�/��8�TKհTKհT��9UKհ$K°F��yA>ˉ/r�)^�]u����`i���E~��X��,A���_R�%X���X���X��E���&XR�%XR�E�yx��.`��.�E�/��_�|p��<�#�R�/�͑�X"�%XTT|����F��[�/���L��/�����e�yW��/���_�7��h��"��i��r�~�l�\�_.�/���/r2�F�\����q�~�Y�ܬ_n�/7�k�/�\���U_�7:'\�_��/�����e���r�~�l�"�o>��_�QCn�/��_��VF|��尢
⋼l痛����y�����e���r�~�l�"��o>��_�!ܬ_n�/7뗛��>�/�~�G�"'������EE�y.��[��n�/�Qw�����]�����<��������rKр�E~��d��/��u_�������㋼ �����������,GE_�7�ObY|����@�-�ȣ:��_.��o�Y�n�/�O�Y���r��񿨻�"��s!_ğ�.`��.�E�k��%X�d|����'㋸ꁥXR��X�b|���H�'�<��R�Eu���>

�z`��z`Q��E��,z2���!Ѝ�E����4W��/rX�Z�E�	�+���E����q2���\�_n�/��}_�C�O|���c��]n�o���}/�=�l7��������z�v��E��k�޿]��.�o�������������E��~[>�m��.�o��?̋<=�2���x����ֶ|b� �`��-�ؖOl�l7�������z���F~�n�l�&�Mۦ��x�G�)m
��`�G��ؖOl%<�q��[v��x�ϔ{ߨW�z�-(x�����l��Vl���
lK�%ے��1��-غ���<�l�l�l���a��%[*��/��3�lA�lA�l���
l^�!�L��m�Ë<�3GP��[�u[�-f�"�-x����l�l���a��]ۮ�mWö�a��-[*������R�-�v5l���>�	
��`
�%ے�-;x��wb���	[���	[���	[���	[���	��xTǶ�-;��>l���l���l��lA���aۯ��[=��[=��[*���o���a�ʅ-غ��ؖ)l����	ۍ�m�¶La��e
[*���2�q.;�T`K�T`K�T`K�.`[��E ۍ�m��l�v���]�߮�o�����/�>�޿]�߮�o�����j�����<�?<E /�\+���
lk�.`��.�E~�SN�-@� l�.`��`� ��E^�#M��������l]��l]�l���`� ���7����l�v��v���߶l�l^�!|$l�l��.`���ۍ����v��E|����Z7���[�E ۍ����v��v����Vl����j�-�n�o7�_�7���.�v��˿�1x��pʹ��1x������E [�]�߮�o�^�Q���Vl�������z�v�[m�]�߮�o���������.�v��v�"�dr��E~���]��.�� a�޿�����ow�����]�m����`[m��6�"�-�"�-�n�o{�`� �`�˿]�?~�x�\�߮�o����/�N8u[��6�R�m����`�v��[*��6�6l���
lK�[=�".[=�m(x����C8}e�j��D�J�m����`�^�Q���m��V5l	Ö0l	��+l��^a��=[���	[���	[��"��+l��V"l%�lA���`�Sv�--�6l%<�s5���l���aK��[հU�V���N9�Ë��>j��ak���E��h�VHl9��>l
^�7:E�҂���:�-��r�]�4���a��a��a���a�^�!V尒Cl9ĖCl9Ķ�`k��a�=��/���l���a���aK��aK����m���{`�!�b�=�[!��#�r�m��VHl9��>l��:l�öU`k�Eۢ����r��}�B�qUöU`��a���a���a���a���a�^���'��[���[���1�6l�ö��E�髐��l�Ķ�`�(^乜�
��>ZZ�u[G��6x�7�gL���b�c�"����d��s9��[m�u/����`l�� c�(^�7:j�[!��[�"N��ت�m¶ a��a���[հU�N�=�4;��a���a��5	ۚ��}ت�-a��-a��m¶ a[���/�\N&�ö a[��[�-@�
�ysCv"l�Ķ�`+$^��&
�m��Ml��Ml���b�(��b�(��b�(^�|�Vliű �($^���Gq�D8
�c'�M���>���bX9đC9đC9ċ<#�XmpǶ�#�8 ��Q�GmqtGGqtGGqtGGq,S8:���8�$��QH���3�QH9ċ� ��QH9đCU�Q5U�Q5��od��ñ��h���b�c1�QH��QH��B�($�����c}ñ��H+^�����E~��Ϯ����^��P��"���iM��d��s9�o82�#�86:��G�q�G�q�/�>1�s1Ǒi��C8eG�qd/�NL{���9�r��4�����#�x��Is����"��೾�(7�r�(7��G�qdG�q4G�q4G�q4ǒ�q.�Ʊ��(7�L�h2�&�0����(����(�h�&�h�&�h�($�B��!����pGq�o8
�c�ñ��E�����8j�c��`K� �0� �X�p4G�q,y8�#�8�#�8�7��o����7�Ʊ��0� �X�p,f82�c1Ë��B��Qn��Qn��Qn����9^�����;^���8F�Ǒ|�Ǒ|� ���X�"�8jm�8Z�#9*��9�>a��aȱ��hE�V�C^�Q�Z�c���a����w}ǋ�l'��G�q�G�q�G�q,y8b����9�}8��#�8��#�8VA�Ǳ
�E�J��Q�ȑ|� �
�@���H>�%G�"�kaȋ���� �0�@�
���pT Grl�8���WN�q$/��r�C��ъ��ъa��a�Q��Q��Ǳ��H>�%ǒ�#9#9#9�CK�
�X�p�!Gr$G�q$G�q�j8v5+��G�q�/⨒��qn�0�C�0�C�0�C�0�C�
�H>���E~��I�q$�F��9*��9*�c���a���'��iZ�#9�9�<a�Q��Ǒ|�Ǳ��@���Ef��Q��0�C�0��;����;����;���9���Xq��8b��d�5����8����8ʍ#�8��qA�,�i�Ƒi�Ƒi�ƑiMƋ�ӖiM�`k%�&�h2����8j���8�C�`ƑViőV��{��`{��G�q4G�q4G��"�H�d��Q[#����(^�Q}��ViőViűC�-���&�h��q�Gq�G�p��އ�j86:Uñ��X�p�ǒ�#t8B�#t86:�Ȼ��PH���>���>��s9M�/���/��,�8��#�8F��M�ı0��(����(����q�GZqtGGqt/�>Y�&�B�($���Z���x���_�Ҋc��Q[��Q[�&� �0� ��(�MGZq��Z���8j���8:�cađViőVi�M��M���>��:��:{����������q�
G�p�	G�p��އ�D8J��D8J�yW|�#N8vH���+�!���H�^��8�Xq��8�#a8�C	ñ
���G�p�/�N�U�*�cı
�EUGqt���8:�cađV��Qű�&��GGqg|�M�ċ<������8j�yTg� �0���E�gL�ű|�0^���:M��dMƱ���4�L��4�&�h2��/�N_1Ǳ��;��G�q,�8*�yTN�!Gr�!Gr�!Gr$/�\Nr�Q��Ǒ|{2�=Ǟ�+�*�kO��\a�U�\�U�\K1^�!�W+r�"W+rU WrU WrU W�"/�}�!Wr�/�L�y��s�jE�V�jE�V��cb^{2�
�@�
�Z�q�1D_�`�^���\a��\a�U�\�.�0�
C�?��Պ\aȕ|��od~]�Ǖ|\{2���J>��׺�+�b�+�xߨ�Vg\�3���ꌫ�����2�+Ӹ�i\��Un\�Ƶ`�E�h�����;���9���9�eW�q��f�+�2�k��Un\��Un\�ƕi\M��d\M��d\6�L�.�=/�Vʍ�ܸVg\M��d\M��d\M��d\M��d\�3� �
0^���(�WZq�WZq�WGq-��Y\�,�h�*$�B�*$��ZqW!qW!q퐸����棏h�*$�B�
�MW�pUw;:$�Z��jx��P�>\U�U5\	Õ0\�&����4�"�*�Tw-��r�+��ڇ+tx���iH�p-��ڇ�}�ڇ�}�B�+t�B�+t�B��j���+a��k��+\���������ZQ�"o��>J�+(���+(���+(���+���6M\A�\A��i�Z+q�����+;����1�6M\���<�S�Z�k��U"�ȏw~)���� ����*��z���F��� ���އqst׍����u��E|�h�õ���mt���_���[�ו����u���ݿ��0\��;�/�O��ԺFmN�n�_7믛�����f�u���Yݬ���	�e�y.��n1�u%��lma��0\W�+�/�}�_�گp]���]u����]ܿ.�_��+�ו��J�u%���]ɿ�俈?m����������uq���]ɿ��_W�+�������u���ݿ���_��_�Q}�q��Z�pݿ�.�_+�������f��_�گpݿ����s���ݬ��+\���
������u���lmN�.ۿ�s9�,S���_��+��~����<��-�kõ��E������uK�گpݿ�.�_�������ug��3�1���_����j���u���Yݬ���_K��/�|�r]�E~�s�u�k���B���"��9��	�����k����F]���ѿ�C8ܙ�n�_���ע����ug�Z4�M���1�����u��E������u���=p��v��s9`�#���_�^�!|�r�������V\���������z�u�����6���_���������z�u����]����O��_�7�����uq����"��uq���]ܿ.�_;����]����uq���]ܿ.�_������5���uA�ZGp]��.ȿ�s��".�}�{��=pݙ���_w����m�k��uA�����\�� ם��>Y�#����f�ug��3ݙ��̿ȏw�pm���__�ݬ����E�{��k��5���u���F]���ѿ�;��q���F]������F}��m�P�3�����u���p]��B>�S�e���u���l]��.�_�����e��f�u��E�ˆ��f�ug�� ��n�_�����V�k��uA�� ]��n�_W�_�!�_�_�ܯK�ץ��R�u]���~�M�.�_��_�_ �����_w�_乜r��_�կ���u���u]����"O�b�կ���E��"�u���~m(�6\�կ��/����������~�`w��҂�~|��n���a�A��0�MK^�{��u�p]=\W���u�p]�E�)�����y�b���+��y�b���>yX4��s1�}�p�<�����h�E^#-\1W�_�V/�\̯p=\D��í� �#�^乘_�zXZn����{������{XZ��{�a�A��{��{�c{�a�A�v����C8��1x���xtA>\�W����p�=�s���=�p�=����u�p]=,7���y|/���[�/�x${��/w����p�<\1W���p��E��i��y�u���+����í�p�<���v��E���s�[��y�b��?|�����?\D���p�<\���M�pS<|�~�<.����ߥ���+����í�p�<|�~���"����	7���p��k:7��>Y����?�s��÷������{����?\}_������7��M�p-<\w���>�ȏw��)��>��l��|��>y�<.������x�������x�)n���5��><�)���k��{�õ�p-<\��3����ȿ&w����y'��?�/���õ�p-<|�|����������y�?��5������u�p]=\W���u�p]=\W�F�����E�p���[F����#?�_'.�:������z��������ῥf#᰺��Ӑ/���UK#���rg>ܙ���p�=�`��R�� '���_n�������h�7:s�3��l�R{��.��K��R{����������oOD���+��y�b��P3��0��=�'�ӌ�x���}�p�<�'�����py<|y{���p-���F~�C�M�pS<\w��w���C���x�)��=\��õ�p<|{����w���p�;\��Å�p�;\���.|G�ԑ�	_��r����;��w����ﯗ����r�oDW��U�p�;\�W�����{��K��U�p�;|Iz���$=|Iz���p<�_���E~�Ɨ��oDW���p�<|Iz�un��+�/��W����py<�7��M�y� �p�;�������p�;\�W��������bu���pe:܏�����p?:|#z�2�L����~t��G����~t���<|ey��n>��,���Pp?:\����e�p:\����e�p:\����e�p:\�~���_:n>����+��e����+�Õ�������_�Q}\���+�Í�p#;��~�Gu~����<���O�m�{���v��.i�K����������v����<��w����������_�Q���_�����u���y.��\�7�Í�p�:\�ׯ�ן��/�N81}#z���_����u�EnQ�[��u�E��<\��O.V�������-�pe:܏�������G����2t���p?:܏��×������_�7���u������;�r�:|?y��nd���Fv����<\����%������Í�p#�E�	��K��v���y<�����׌����k��U�pI;��ׯ���p�:\�ׯ���p�:\�ׯ�]�p�:|5x�~�Z����u�k�Z�+���t��"?މ�K�×~����bu�X�.V����bu�j�������3ݵN������,|��,L������^S.]�~�ϳ\���nd���Fv���nd�/�N���%�tI�E���.i�K�����W�����Fv�~��_����������t�:}�w�X�nQ����2t���n>�k�鋺�5�y&S����4���Nw�ӝ�t�9}ww���"?�㋺�u����r�����;�VN�ݝ.0�r�,����y���v�����;}+w�V�t��E�q8`�|~�w�i�s���t�9}�v���"�CM���"?���+�ӝ�y����/�\<��/�~��r2�X�.V�[��u�E�"��r�:}ww�X�"��]�t�:}�w�k���;]�N_��"/�a��u���t#;��N7�Ӎ�yz~,�{���ӽ���/��XL�)��@<]�N_ �;�/�~9�\O��ӵ�����x��.|��/��+Y�ݝnw����*w���.i�K����_�!���m�{���v�����<]�N�O���<}�x�ݝnw������ӗ��/#�w�g9_3�"�8�'O���}��5�/��u�n��+��>���x��+��>���xg��'OW���y��.�����"��<��w��������yT'���{�b�t�=�`O���u��-��[�ӥ��-��R{�Ԟ���E���R{���t��E�ˉ�6|�����q<����������{������K��R���Fg���/���MOw�_�Q]DO�_�g9�S���N��s�=}�z�������s9]���x��Bw�ӝ�t�=�sO��_��;�\jO��ӥ�t�=]jO���K��R{�Ԟn����+��W���xO_ޞ��=]}��p~� ���=ݙOw�ӝ����+�����K�/���eO7���t�=�`O���.��/\O_���p=݆OW�ӷ��oWO���yT痯eO7��������}�l�.ۧ�����_�Qi���sO���e�����k�_���{'|n�[��~����=]�OW�ӕ�t�>ݿO���"�S����ȣ:���Ow��]�t�?��.����]�t�?]�O����tq?}S{�����=}-��8W�x'H@�>�t�?]�O���"�8|�{�������N�z�E�ˉ)H�@Jҍ��Y�/@�>�yz��. ��O7�3�_�����H]@�R�"��,Lg�z �/��B�@���T�z ����ӷѧz �/�O����/�3��g�]�7�����Wϧ!}�|�^�7�R�T"�o���ȝ�=��{���̧o�O� �ڇ�>��!}�|���y.��"}�|J+RZ�:��Q��"}�|�(RG�"o�CT4��T>}�|����Q�������Q�h"E�K�SG���TH�B"��H�D*$R!�r�y.���7ȿ�s�SWZ�Ҋ�V��"�/��diE�(R4�"?އ@9D�!R���>��}H�C����C�"�)�H9D�!�7ۧ"���_�|T�5��k�ӷѧ�"u��H�D�&R4�"/����SZ�:��e�)�H�l�ҊTH�B"��H_v����e����ӗݧ�"}�}
0^乜���L#5�Ϗw�	0�7ۧ&#��S����`���O�E�-R4�
�������r~��J4�"�N�(R4���M�"��}H�CjRՐ�z>����_�7:�|�|
^�7�o|B�:��!�)tH�C���y�_��>�)tH�C
R�B�:���E�{�҄)tx���)�Wϧ�!�)tH_*��A>�)�H� �"��H��}(�C	J�PB�:���|���~/�E~#S���}(�C	J��"����/���C��|A}�6��C���%�(�C	J�P��_%N(q��̯�+�?���WϿ�C�U�z��%t�̯�=��{���̗�|�|)$J!Q
����%�(�3_����(E���V�o�/�E�-JmQj���(�EI+JZQ�.����(� _�A�|�|���i�&�|�|i2J�Q����/��B�Fi2�WϗL�4��(F	0J�Q�g����(_=_�g��/�:���ԗ/�/1G�9J��"�Ĕ|���/H�@JR*�R��
�T �)ȋ<*υ%�(�GI>J�Q�K�T �)H�.��|��Clǣ��E�q�.��|�䣶�QR���T �)H�@J�Q���w������(߸_2�`�ڢ�%�(iE�(��뗴�|�~�-JmQj�R[�ڢ�%�(E�J���%�(iEI+JZQҊ�-���(iE����V���/ŋ�F痴��%�(_�_Ҋy��j�x'�(�ŋ8�h�D�{�_��;��nҊ�U�%�(iE���񧭶(iE�(JGQ:��Q�h�D%�(�D)$^�����;�KQ�п��x}}��&J4Q��M�h�l(E�(����B���(�D�!JQ6��l(�DiJ�Pڇ�>����㔳	��;��w����/E�(�w�����/�~I+�&��	�E�)'�(iŋ�F����t��(�JQr���>��*P�
��%�(iEI+JZQҊyT'�E%�(EYP��M�u��(JGQ��M��k������(�D)$J!QV��l(�D�*PV�uX�&J4Q6���
g�ڢ���xw5|Jǐ ����(�E�=Pj��V�B�/����3�D�&J!Q
��C���%�(9DYG�"�M�h�%�x��胛B��1({^�pX)$�҂M�h�D%�(�D)$J�"�H�C��C8���(�D)$�j�RH���e�AiJ��">+�r���ڠ�a�j(UCI^��R5����D(UCىP����T�j(��ys�_r��>�%�(9D�vPڇy��/J!Q
�RH����j(J�PV�8�E~�?m;(�B���yW}�� �T/�:���}(�CiJ�Pڇ�r���}(�CY�P3�-%�(9DY�P
�RH�B��e�Ë<��wr��C���%�(�C	J�PB�yǣ�%t(UË�F'����e�D�!JQ�J�B�E�Q��(�'J4Q6M�h�D%�(�DY+Q��y'����M���E^�CT�P��0����
%N(qB��Pz����lt(	C��P��R5��/�F�^�!�e�CiJ�Pڇ�>���T�jx��p�J�P���
�E���}(�C�!Qr��C���e�D)$J!Qr��>���E���v�Y+Qr��C�Me�D�&J!Q
�RH�B�%�(�Ë����T�PB�y�Q�(�>��C��,�(�CiJ��ƪ�p�����\�����(E�(�l���(+*JmQj����%�(�D�&J4Q�J����(E�(�v���E~�SNGQ:��q�#MZQ���0�t��(E�&�*�M�B��a5N&�ċ��+iEI+JGQ:��Q��%�(iEI+JGQ:��Q���t��(ŋ<�SNGQ:��Q���,�(iEY>Q6M�ڢu-�x��߉M�h�-�x��5�-�x��~#O|-�hiEK+ZG�:��Q��o�_[+�"/���Ҋ�V����m�D�-ڦ�`�Mm�D[+�vH�r�E����i�L�e-�hMFk2�>��i�L�e-�h+*Z��2��i�&�5��hMƋ<��/�ǖi� ����h�,Zm�j�q�v[� ���hiE�(^�eK+ZZ�6`���E-�h�-ZG�:��Q�u-�x���[N9iE[w�j�����-�hiEK+�n����E&�hE�(^�e��j��V������rҊ�Q���u/�\<����-�hiEK+�΍�s�-�hF�-Zm�Ҋ�V����h�4Zm�j��`��-�hiŋ�xg��-�hiEK+ڂ��`�-�xڶi��C85m�F�4ڂ�Vn�/�Z�3Z��b��'��-�h1ǋ�l����x�M��b����mOF+7Z��ʍ�i�L�e-�h�.ں��i�L�em)Fk2Z�њ���e��hMFۀ��]�&��h�F�4Z�њ��d�/�m�h�F�4Z�іb��s����hMF[dњ��d�&�mEk2Z�њ����5mE�&Z4�r��C��/�9�O��-�hiEK+ZZіO�ڢ���h�E�-^�QiVT�-�h�F�4Z��2��i�L��h�Ƌ<��P��ʍVn�r�e-�x��:���h�3�ꌶ:�E�˟͒��|��-�hH۹�vn�V��"m�FۦѶi����"�i�HkEZ+�"��֊�V��!/�\Nr�H���򑶿��#-��p���|��#mG+JZQҊ�V��e}�� �I����w�:��)-Ei)J[��ꔶ���)/���$��u�kX^��r�_Ƕ%"��i�K�_Z�������5,m�H�ZZ�Ҳ�����"�tiC�Ɛ�1��0��i=L�aZ�z��ô�mi�̋<�9���ô�E�m�HKd���ȴD�E�z��j��i�LKdZ�����!��iCZ"�6��j�U3��i�̋<��7��B�Ҵ�"m�HKdZ"Ӗ��%"/�N8j�imMkk���鳯�"m�H�rZ�Ӣ��۴ܦ�6-�i�M�m^Ľ�W��6��im͋<���r��}�8��i�M[5�B�Ҽ��r��+�B��1�mimMkk�Ɛ�۴�!m�G�fZ5Ӫ�����4-�i!͋��>
iZH��N��j��i�LKdZ"���ȴD�-i�LKdZ"���1�%2mcH�fZ�z������/�ti�J[�т�֝��u'�;i�I�N^�!�AlYG�NZwҖu��u'�;i�:ZQ�6s�Ȥ����1JQҶi�m-2iEI+Jں�V��ț�L�I�L�R�yW0�ѝ����h�I+JZQҊ�V����%�(iEI[��"����-2i�4ZwҺ�֝�|��#��_�̤(iEI+JZ>�򑖏��(i�H�G^���Ƨ(i�HC�ꌖ|��%-�h}G[w�v[�ȏw��;Z������%m�E[w�*�V���%-�h}G[�ђ�s�/�����h}G�;Z�����w�m/�\�/�4Z���d�
�U �iȋ�8�w���iaH�@Z�Ѷi�����h�3Z���yT���m������F��ʍVn�r��m)F�9Z��ʍVn�ȣ��e)F+7Z��"�9�Ƌ�_�/K1Z�����w������h�Fۓ��s��c��1�(7F�12��c�c)�X�1�����|��c$#�1�Xw1ʍ��b���M�h2F�1��`� �E^#�2?Vg����\��d�&c,�6F�1ʍ�ǿl�m#����4�������h2F�1�i�Lcdc��(7F�12��d�&c4/�\���:c����X�1b�Qn�r�E�K�12��i�=��{2F�1�d��c�#�K1F�1��`� c��-F��"/�Y�����4F�16`��ot�)7F�16`�Lc,�M�h2F�1�`�uckŨ-FG1:��Q��bD#����!F�0B��Cb�#t�Ë�l��^�ǹ������($�>�q.+*F!1�O������($F!1ڇ�>���}x���:��a�/��� ��jUè�֊:�}�jU��G1��Q5��C8�l�x��r2iF�0Y�b�#��,F!1
�yz�D#��Ĉ&F1Y�E#������>�}#�9ċ��ڇy�b�#�9�Xd1
���bD#�9ċ�x���L41�V�h�E^���֊9���Q��?�}c�($Ɗ���b���X>1�O��bt���Ĉ&F41��M�hbD#���F�0B�:��a�#t	�HF�0���b�U��41z��+�^a�
c��HF�0��0��a$#NqF�0�����E�	R��"���b�	#Nq�֊Q"�}�1���F=�"O�#��#(A�
FP0�Q�T`��z��41������z���?���}�����?.�[�����l��uX�Z1�ߏ��c�ċ� ��Ǖ�q%\�W�Ǖ�q%\����drK�����-�qK�����-�qK��W��֊q%\������q�~ܬ7��>�q�~,��'�5�q��E~���>�q�~ܬ7�ǝ�q~\}W����q�}\}W��q�}�;$�m�q~\}W����q�&��qA~\���>�qg~ܙw�ǝ�qg~\���rZd1nֿȣ:ݬ���Y���l?�]���cƸ�?6`�+��J��<�Oiv[���/��}p��bܿ���֊q�~ܿ�,^�]ub��?����/��-j��Xw1�]����.���?����J��m1��+�c���m1��Ec�Ÿ�?n�[��J��C�-�qK����-�qK,����-�qK�x��r��"��Y�.�Xd1����;����E�ˑfE�XQ1R��
�T`��]���>��
�T�E���+���c�Ĉ F06M�M#x��rb��Q*�"?�)gE�
FP�"��Qc0����[+FP0�Q����BA�Xd1����`#(x���s�z`��;$���CbD #7��Z���c�Ĉ F0"���s9�D #k%F0�J��#k%^�|��Cb��x���H��;�H�Vbd#;�&Fv0����`��#F=0�Q��/��r����c��(F�0J����`4ca�
FP0�����^��rꁑ
�T�E~��O=06M���vZ1���Cb4�1��X+1�J��`d/�VJ��V�E�	G��a$#a	�HF�0��0��a$#a�Ʀ�'�8a��D%�(F�0J�Q"��`dc��X+1�'�8����W��et��Q%��,�"?���������_�����"��w��w�}��;��;��x�EM�;��o���_�]���_�~g�~���k���_�7���/��y����E��w�}���|_�_�ߑ�E��w�}���|_���|_�~������������<��,�"��;����;�ȣ��/�N9j%���_�n_�Q_��_�-��<�#m9Җ�Z�/�\��_乜�x�/���T�E���D�"���� �E���|�����E��!���F_�~_�,�0|��r�-�_乜�؇/�\���,�|�<��~��w<�&��s91���"��ĤV⋼�NL �yW(���;D_�Q��GE �q. �q.L�qTL�qWa_�Q�t[|���@�d|���o�_���{�I�逸i⋼�N��c�v #7��C��	���?�p #7��������C8�a/rԢ-���C'&���x'&�⋼F����m�"'& �<�C��E�Y���"�,���<����E���Ǚ��"�
��"����"�_�!V8�/�ί�% ��8���JZ+�ȣ:� _�7:�h��"���Ek���>c"7��C8�`_�i�b��gL0�yT�1��x����E^�S�8�h�x����E�����?�ѻ�B[|���w-�"���E�U
#��C 0���`|��r^g!�⋸�C|���g3�_�p�0�ț�H�
�E�{! �<�OiЊ/�N9��y'��L}ËV�_�h�/�V��/�98�/���]K��y��E[|������F��hN�"�d�V|��LЊ/�}��&ዸ4'|WiN�"�
��"΅��"����r�<�#��E�ˑ��x��r��/�Vh�9� _�������d� ��F�_�!|p�i��G2���Y�/LƋ|�
��a���"?����"o�OV0�/�r0�9�`_�Q|ȍ/�>�c�E����"o����E���E|#L��x��q�h�/₠_č�Q���8�/�V��/�_�/�Vp�/�Vp�/�����>YQZ�"�h(�"�c��E�5�u_�5�����t��(^�H�Q|�Gu�!$��s9��1�"?�Ʉ}�"��1��"��}J�>|߈j�">�:�/�O��E�:�9��
_��;��g&�Ë�L��/�N8�P_�V�:|�7��؇/��/������>��E> �c�E��(p��Y�!p������8�EΜ�1���/�\�8��F��
��E~��	��E^��Lx�/�O�ɄW�"�8�_��#��o'|w���E��y���C8�ڑF��y.���<����E�5� �<��
��E�ˑtx��_��/�i�#�ዼF� _�!����/򲝘��/����/�}$C5|��������x�/�:�h;�"?ޑ�W�"O��8ዼF�S��E��/�㔣��E�������H�9��6�"n!��F�����F�QZ�E~�H��/�C��/�Μ�g �<��_�d�+|�Gu!��C���D�"�d�|��r�Љ�E~�Oi��/�V��/��/���V�/��LP�/��V�~\��E����kI�T`I^�{���E�g�Es�y.ܖ�`Q��E���DX��y'�/���%NX�E�����^#��E~<�dK�����/��%NX�%NX�%NX℥DX��%;X��EM�yɖa)�a)�_��3��`i��`i��`i��`i5	_�����I�"��]��E'����HM����	Ò0��o�pI�^�}��[�[�',q¢��xG��`i��`i^�QV��1X��XR��X��/W�������f������FG_�vt�F�\�_��/w�;���Ei�y�?���3�;�˝���rA~� �\�_n�/��_�!� n�/
^����٦{���,jh(�"OϿ3-�^�p�}QG�E�	9�s_�/���t���4|���ߙ�{��=�7�=��^�7��CC�ys|�q�~�F�ܙ_n�/�����m���r��E^��9t|��p�m~�-����C��E_�5�E_Ĺ\�_.�/����E��y��;󋢁���5���r�~�F�\�_��/��k��5�����x��\�_�|���9w�;�˝����rg�E�˟���/
���;1ݙ_.�/����E�y����/w�=_�7��F��y�N9��������F��y�>˹Y��1�"���r�~�3�܆_n�/��u_�� ��#�"���=�E^����E���Y>���h�"O�dr��E�aE�����Z��ot� �\�_n�/��E_�7::\}_����k���:s�#�"�љC����3� �\�_.�/�_�7:��������r�~�F�܆_4|����r�}����s_�/��=_�e����s_�/��_�!|آ����9>Y� �\�_�|��rʹ �\�_nÿ�otʹ �܆�w�YN�p��c�E^�OV��/��k�҂/�}�r�~�l�ܬ_��/w��j��d�6�r�E~�S��E����r.�/��/�>w�_�_ 
�����EN9�_�5RG�E-�^�OJ���C8�\}_��/W�M _���0�Ln�/���C�c1�Ln�/*��[�drA~�*�E��/7뗛��5�E��y.痛�����f�r�~�Y�ܬ_�|�G�Y���y.e�l�h(�"��࣎���8�7�Y��rK���"�ёF��n�/W�+����/��B���ktq���\�_��/W�+��e���r�~�l�\�_.ۿ�C8D�g9W�+��:�9W�!J�����\-���#x�s���E��y�j��W�Zz^俸I�.`��.`��.`��_��qb�S*��6x��P�tK�"�Ĕ
,�����<�υ�s!=_�!�K�D �����(x��X���x��sa;��_n�/7����������rqQG�E~�#��]KC�y�>��_��h���[��-���rK�����_�|��p~�����_��/W�E_�7:��x��r�
|���dj'�������z�r��޿\�_�|�GuXQG�E�?4]��,����Eίq~� ^�5��`�=�E~��I�\�_��ȣ���z��h�EN&��_�Q0.�/���[�˕��J��<��Q.�/Z^�dr��˿��_��/Z������z��U�E�������]����rqQ!�E^�󋾀/�_��,���s9����n�oW�+�ە��J�v%�E�׸���n�o���[�ە��J�v%[�"��vq���"?�)�]���l�����e��f�����5������l&�v��E�	1���������v��?[w��ƮcpKN� ��o��TQ=�����l�T��ղ��藌~�藌~"��Y��/����~�藌~i�@~��~��~�˿�K �>}&���藌~�藌~"���_~���"��d��/�� ��KY���_2�%�_v�/;���~���~"��_���k���~"��Sڲ�I�$I�'����Y(�_V�O��;�l�_��/������U���rU`�*���_V�/
�˅��B�r�`�P�\(Xn,�����e��r�`�P�,�_�,w�;��e	�r�`�c�\(X6�/���˅�e��D��&�Nظ�lܟ�+���r²�����DXV�/7�%����¼_�����r�`�c��1X��/���;�z����zh>����U����q�=�l�_6�O�p�v��1X.,
����eq��"_��dK�r�`�v�\;X�,w���qE
��U��^�r/`��\X��%�_��%�_ေ�~���_���|��+�K y.��§4��{�%���r	`�����J�%�_���|�+y���/y�D�ɤ�_��%�_�/��'�>���ן�s9��X6�/
�˅��B�r�`�P�\(X.L�Q���/w�;˪����������DXn"L�|psa����DX۹j/����˿��_��/��+����r_aYտ\aXV�/��+�}�eU�D¹j��r�a�հ�WX�+,����
���e{�r�a����DXn",7������B�r�`�P�\(X�
,K����U�e���q٥���_v�/w�;˅�e��rU`"_��/� �K K��_.,� �K �%�%��C8'�y�{˽���r	`ْ��_��/��R�/I���/I���/��$I�$Yc��_v�/I�D�G�sT�K��_����_����_����_v�/��*?͕�f�e����~����	��pYv���K˿l�_��%�_���<���������9a%�r	`"���r/`�0��r~�=��Xn,���yT}l�_n,����큉|y���~�Y���Kl?�??͉헌~����KF�d�KF�d�KF�l����谲�~i�e�KF��_�u�Ԥ��ȗ�9��e���O�0�/���/���O��;��K����K��l�_j���_j���_j��<��C ���K�t�����s_:���>lIߗ�}Iߗ�}Iߗ�}Y����K����K��,�_�O��r�i�f~i�~ْ���K���K���|:�%j_
��`_
��`_v�/;뗂}��'��}��~�Y���紏>:��s_��/����/��ҹ/Q���/��'�C
��M�ȣ:s�_
��`_
�e���/���}�ܗ�}"�ꓕ�}�Y?�Gu2�l���K����K�>��pIߗ�}iӗ6}YP?7Z������_��%j_���`_6�O�}�R�O�-�/����y����J���K���K��_�e��D��/���/����~��@~��~Iߗ�}�ڗ�}�ڗ�}�ڗ5���%}_:�����I���K�>�o�a%}_��%}_��e��R�/5�������°?��e}�b��̇>��;�C j�PÇ��!��|��f���>��}��'�|be}��������C����߇e����<3��a%~��C�������?,��(�'��<v����@إ����O��3}'�<��?l��}(�CY��Pև�>d�!�}��Â���>,��C��ۇ�>��a�}(�C �8��7��O��L�؇�>l�e}(�'�\<���>d�yEǐ�>d�a�}�C ?����y$�|�'�=:�`�D�/>,���!j{��C���Ц�6=��!D�yXc?�/���<$�ag},}��!�x�lJ�P��5�y��rN,>ͅ5��'�xXP����x<�;�Cb󐘇��ag�D��ib�}�Y�󐘇�<$�!1�y��CO���&��P���<,���D�1$1�yH�����O��V����a�}�ò�Ц�6=,���'�4���f�P���=�Q{�Fr����\}"_�)'W;�C�r����\=l�{��C�r���>l���r��]^�)�`{(�C���G���BQ{��C�r����!D�y��Cb󐘇�<��'�Cb��v<��Cu>�R���<T�!1�y��Г�5��'Yx��ò��������x(�C)��L��)��x(�C)���>��a�}�z�<��Ob�O�}��%"�蔳8?,��z��'�\��G��,Թ��=t�a�}��C���ЦO�]��>$�!1k��������Mmzh��6�P���<,��ȗw��Cu�󐘇�<ҙ�:��C�B���=��a}X=r��g>�a��D^�i�`��D�!�D:'t�s��������=D�!j{���P���=��!Wmz�Cu��P�O��T>��qT��Cb�Г��<��!�x���R����!�9��|��;�ݡ�)�D^���w�'�=����ú��~"���a�{��Cb󐘇�<��yED�s!z�C�>���\=��!W�zh�Ê����\=��a7|�vÇ�=t�qT��ú�й��=��{X�Ň@>�!�K�C �ʇf>4�y.���>d�a�|X*�ȇ�=t�a�{���8���!Wk�C�r�Ц���*�ГO��kyT��x<��!�x��C<��p=,\��d����:��+:��GK�'�J����P���|"�W;T�a�z�C�V��%�aIzH�Cb�Г��<��'�x؈>�w�'+��D�'���J�>�7�ǨvY�r�Ц��<T�:�y��Cb󐘇�<ڙc�zX���P��R<�M�x؈��=lD�Cu֟��<T�:���^}��!D!�D�G��C�V��U�Mmz�Cu����<$���4�yH�Cb��<�3GV��U���Ò�P��R<lD�x(�C)J�<��Qz�ГO�Q�q����<�[����<4�!�uwH���{K���{��[���[ʽ-Iߖ�o��D���e�y���|[��e�[�5�[��[�=���ak����[�5�[�5�y.�ז�oY���O�xJ�J��J�-߲��޺��޺��޺�my�io�۷n{�'�L�-��R�m��VwO����|okٷ���Z���ֲo���o��V�o;طx|+ŷ��[���[ݽ��[ݽ?G����v��|�N9�շ��[<���[)�mW���-߲�m��V�o��V�o;ط�[<������-���-��+�,���yG�M�[����[��-o�B��:ߪ�m���]}ۮ�%����|C|��C�Yt�շ��[��-\��-1�v�o����o����|[l�m1���#D�B�m����|�շ\}�u���y.'�\}�շ��[���:�
���9N&Q��}+ط6}kӷ}�η�|�η��ۮ�m��V�o�η�|K̷��yEj�����-�V�o=��o����|�ɷ�|�ɷ�|�ɷ�|[Y�e�[���[ʽ�,�V�o��|O�rN�5V�o+�'���|o+˷|k��|����{���n{�'��}6��|[F���[����N�-��"�-��"�-��6�O����Dʽ������6�o��|o���f|k��|�)���[ʽ��[��u�[��m�R�-垈s����{붷n{[����qE��[����+:Ҭ������߶�oY���oY�D�Y��J����B��|o��|O�p<n�t�[���[��-���;�t�y.��{K���{"O�#�v�YY��S��-��C��(��V�o����|�b��,���-�ȗ�3��|"�,��o��D�g9ѷ��ۮ�m���o!�D^�)�:�v�o!��o!�V�o��D�_=��'�9������!�W�$���7}"���|K̷%�[O>���r)ŷ]�ۮ�-���-�֟o=���|�ɷ]�[b�%�[O>wUb��:��I�N&�η��yEg�6}kӷ-�[b�%��~�m���o�Ƿ��[����[�>�w�#W�r�m�V�o���O���1d��O�pi�'�N�YT�>��w~�ܷ�}[��E�[ԾE�y���}+ط�}�շ6}kӷ6}ۛ���[u���[O���[<���[<��R�V�o=�֓o���o���o�ԷR|+ŷR|"��/�,\߲�m��D���O)�-Iߖ�o�Ϸ���b�����hg�|[Y>�o��ae���|[Y�%���-1�V�o+˷�|K̷�|K̷�|K̷�|K̷�|[Y���[<��'�z���۶�|"�v;sl1���-D�B�-Dߪ�:ߪ�:�󉼢�b�m����g~��'0����o=���|">�-1��-1��-1�z�<��Q��-1��s��dI��oKҷ%�[����[����[����yE��]��b�`����M�B�m���o!�V�o��V�o�η��[�e��~�m?��o���O��o����|�O����2�|C>��·e�[)���[)�-#ߖ�o=�D�	���|_'�e�[��U��2�m�V�o��D^�ce��o���o���@|[ �-��s��b[�V�o���R|+�'��)OYx�����T��R<��O��D��J�T���O�x*�S����CMZ���Ԁ��;�ݩ�NuwJ�SʝR��;��)�N)w�S���y�u�i�wZ��y��;�)�N�wZԝ�|�?>ͥn;E��Z|NK[�'�1�&���g"���S��|��{"޶��)�N�w
�S𝶅�<mO��Ӷ���m�i[x��SO�z�ԓ�m�'O��D��R)�J�f<��)O�x�<�z�ԓ��<��)O�x*�S)>����,��)�ț�Ĵ�|"��[��SO�z�ԓ��<���ȗ��-��)O�x�b�����<%�)1O�xZl���T��]�i�y�u���(1O��D��r
���ԓO���'�|J����<%�i�y.'�]�)O�x��S<���+��D��g9=y�u�v��-��ȣ:M��ieyZY�z�<5�i�x��s��O�xZF���<�OV��<��'O=�D�9>Y�����y<��i�xJ�Sb��@<U�)1O�y���-<��'O�S)���g���O��Ӷ�ԓ�x|"���J8:��'O�x*��:���x<��)�N�w�ݝ�ԀO��#OYx��S���r�u�)�N)w�ʝ��Tw��;�ܩ�N+�S��Vp��{"~���Tw��;��)�ȣ:M�ݩ�N)w�S����_��z"画C~���_�E�yT?"�S�����m�n;u۩�N��SʝR��{"O�Ӑu�)OYx
�Sݝ��i�H{"o�5�?�촨;�)�N�uʯS~��s�"{"�D:�D�ix��S����_��:U��0�y��:-�N}t�S��贕;��N1�D^�ib+w�ʝ*�<�Fk�Z��Z��:�֩�N�'�>3ɯS~����;��i�w���yO����I��6|�n{"߶�L�촻{"�3G����TdOčVd�";٩�N��D^��(����;��)�N��Sk=��w2��p�_��:��)�N�uj�'��/K�SE��~�uީ�NuJ�S�b��4�E�)MNirJ��V;m�NMsj��V;eΩiN��Ӿ�\;e�i�vZ��b�T>O�!��)sNk�S�2�6;�ϩ|N��B�T>��9��)sN�sڑ�2�9���i!v��'��;s�͞�]�\Μ�ӐM�)�N��D��3�8s�֩�N+��
�_��z"���![�'���E�)�NauZ�Z��Z��:��)�N���r�|��㰒L�d:%�)���{����s	�SX��~��:��i�wj�'�N9Ev*�S�����H;E�)�N��'�����MʝR�f|"�S��r���m�m�)�N)w��S�����n;E�)�N�v��S�����H;E�)�N��D����!*�N�vZ ����m�5��N�vZ3>���!�}|�e�)��ț�|��;��i�xZ3�֌�5�i�x*�S��TwO�k9��i5xj�Ӷ𔅧,|"��H���O�xj�S�=�/���~~TwO���e�x
�Ӛ�Ԁ�<5�i�x
�S�v����Ox�������ix��S��|"�Ŝ(uw��K�]���m�n�tۥ�.Ev��]�����C.��˾�_�ֺ�֥�.�uY�]Z�V����ե�.�KE]*�RQ�d�$�emv��K2]��L�d�$�eGvّ]b�����e�u��'���Pb�?���d�$�%�.�tI��B�RQ����ѥ�.}t)�K�\��R>���yg�̹l�.�s٤]6i��l�.1t}�!�sɜK�<�Wt2i�����4�Z���.�r��K�\V]�UץV.�r����겞�>J�\:��	��ƥ0.�qYO]r�����.�q)�Ka\
�8��x"�C.r�K�<�&��ץV.�'��;�K�\���4���,�.s	�K�\j�R+O�{t樕����z"_�O:%M.��˪��x-���׺�ʥV.��D��˪뉼��9��R>��ϥ|.�sɜK�\�f��d�y'�L2�9�̹,�.M�D��̹4���y"�j8��ϥ|.˵K�\2�\�,מ�s9�nVp���$�ewY�]Vp�d��ѥ�.}t�˾�|��W��<���l�.uY�=���)�r�b+�ui��7>�e+wɯK~]��_���Tԥ�~��i�V�f�oB4�=:��a��.Ev)�K�]��\��e�v)��#y��H�D�%�.�v��K�]Vp�n�D�%�.�vY���:�ț$(uw��˾�|����.x	�K�]R��m�H�Dڥ�.�ui�Kk]��W�h�i��W�g��_Z�#���%�.K����W�b�p�(�_��W�G�>��ѯY��9��.}tYO����"�9a�uɯK~���<�����f�"���e=u)���'��EZ�RQ���Џ���1t���#���e�t)�K�\��9�����r#_�'���겞���.�tI�K2]���G���ￔq��	�z��G����.}tYO]�S�����EF�8�e�Z�H�Dڥ�.Ev)���9#��G7Ev)�K�]�����e�u�~]V]�Uץ�~s�����4�v��K�]�X�n�,����G�s���l�.�K^��Rw���t�e=uI��z�r��{"߶�'�ĺ�%�.�w	�K�]�_���e��D\Q^�Ҁ��4�e�uYu]��|�໬�.xi�K>���~9��/�x)������x���/˵'�>����%/Yx��K>��7���l�.Yx٤]J�R��R���%�.�w	�K�]�k���e�v٤]�����ڥ'/��Kb^��8�����'/=y��K<^����x���/�x)�K)^J�R��,�d�/x	�K�]��|yG��%/K������x���e5x��K<^6|�x���%/�x��K<^��R��uޥ/�x)�K)^��λ��.�x	�K�=�r�G'���tۥ۞�B�#�}��m�n�,�.)w)�'��!�.�'�R���,�.�w	�����{"O���x�l/=y��K<^��Ҁ��,/�K)^J�R����%/��񒘗�:/�yI�Kb^�S�T�:/��D�/g�5�:/�y�)^��R�O�O��ב�'/��˚�<��O�^B������%D?B�#D?��'�����Ѧm��S|"��H;���<=#��<~l?6���'�<�M�Q�rGF4�G3�,?2��<O|GY�,?�x�;��#�?2�#�?2���?��#��ȗgkƏf�h�f�h�'�\L�#����_���c�������kƏ5�GY��y�厲�(�@��@�X~�G ���>:��s?:��s?�~��D���G�~�?��{������X�},�>��c����O�CV�K�����菥���?����?2�c�������'�<F����O�!i[G���:�c����O�v~}�/���O��Hy��GY��GY��GY��g9���K��Gl��Gl����iˑf[�D�{G���X ~��G�?2�c�������'�9�l?��c[�������~"�3G���0����?����?b��<�H���<��Il��Gl,?���Q�O�ˋ폝�q��������������X3~��Gl��GYl?��#�?��e�Q���'�F;����~�#�?b�#�?b�c?���������D����yE����G?�Wt�I���G�$�y~Y��G�T�ǒ�#�?6�-���O�|��Kҏ�����v���������؈>��p�)돲�h�@�l��@���'�N&5�Q�5�Q�5�Q�5�Q�5��������XY>�/ϯΏf��b~�,?2�#�?2�c?�����'�\~�S�e���[̏-��������b~l1��+�i�b�#�?v���Q�[̏-�G���G�$��-6��C8���G�T�G���Ǯ�?�R:����F���?֟�Ϗ�~">֟�Ϗ$�H�]�G�,6?����������D�{}l1?��I��l1?����Q�����O��vX�p��qEN&��Q��͏��G��,?*���?��ce�Q���Q�O�!0*���?����?��cI���I�������h���b~l1?����~����h�f~"��D �yE��f�h�'�~���O�p�X�~�R?����?���<�CA�~�G�~�,�������|"~B
�#W?r�ce�Q�[̏-�G�~��G�~��G�~�,?�#1�ȗ������Ώ���ɏe��2�#?6��Ǐ�|�?��O��a���y|"�?w������S��)~��G)~����><(ŏR�(ŏR�(ŏ��G~4�G~��G�=oH�}D�G~}��G~}l�>��c�D��iE���{"ᜐ_���Za�D��CAk},�>��#�>�꣢>��c��QQ;�������W�I�r�#�>6i����z"�地6�X�}�����#�>��/��D�Q�&�#�>"�#�>"�cm��_a�V��L���L}��G}��G���d�H��d�ط}��>��#�>��#�>��#�>*�s�_��#�>��#�>��#�>�ꉼ_��F~=��w<*����ȯ���X�}��G~}��y}�i��DՁl��D��[�!z��퉼�CT�}t�G�}t�y.���{"��xl�w[3���Vw�����-�n)wK�[��R�r�n�uۭ�n�v�[��"��u�����R��m�n�u�ys�-�n)wK�'�\�ǖr�?�D�<���-��ȷ�,l�w[���Vw�����mIz�ے�ր��5�-�n��D^�Y8��`��5�m�z�[�݂�J}"���c��[޲𖅷,�5�mozۛ������y.�1[b�󖘷ļ�Ro�yK�[O����R�����_J�V���5��n�v�ۮ�VdO�]�ɪ�֭�n��'��|�N��g���&"�$�E�-�n�uk�[kݖ��%�m�y[�"�i�H�E�-�n�v��[�=���aK�݊�Vd���-6oEvk�[k�Z��Z�ֺ�?o�u[l޶�O�}�i�H���m�y[l>�?Z>��ֺ��-��圐L�d�m1o�tK����L�d�%�my/'���Vn�r����0��y"~�����5ͭinMsk�[�<���@��v����-sn�[����V>��y"���C�� �n1t�<���9���5ͭinMsk�'�m�I�<�G�#�e�my˜[��2�0����-`ns��'�F�#`n��D�a%`nk�ۚ�f��oMs�)ޚ�0���m5x[��0���m�wK�'��r���:�V+�Zy"���4���5ͭinM�D�O'�y����-`ns[��vw���yz#�0n��[t<�G�����mww��'���}��FD��:��=�y�X#:n�q��[t�������-'n9qˉ۶𶻻���?�-T�u�-:n�q+�[N�vw�¸�m�w+�'��qˉ[N�r�����ín�pk�[(�B�
�Px"��4�����ín��[N�r���x"��̑���0n9q[ �
���o��D�|�qKt�V���E��E�-:n��[tܢ��u�m5xK�[��:��!�踭�n�'�V��&�4�����#�u�-`nirK��:�λ��nir�'��V:���ƭ0n��:��{"�c�:�<��I��涨�5�mQw˜ۢ�9���-�n�s˜���V>�u�-�n+�[���m�Z�m�nirۑ�vd����-`ns��8`��n�D^љ#snk�[��6iO�p�h����9��y"��d�o{"��2+��
�VQ�d�%�y.��d���nu��'��/u��[2�6i�d�mҞ�+
����xyau��ێ���Z��Z��-�nEv+�[�݊�Vd�"���-�n�uk�ێ�#���n�v��[��Z��ZO��k��vX)�[�=�o�O��k��n�u�m�u�~ݶ_����ܭ�n�v��۪�i��׭�n�v�[�ݺ�i�H���n�v�[~��� ?��/�D�m�vۤ�R�6���-�n�v+�[�=���Rd��z"����!u�Eݒ�L�>�e�-sn�s˜[��VJ�����}j�V+�Z��ʭVnirK��:M��>VJ�Z����oϗw��[���0�]ԭinM�D��ins�X}��4tm����~�x���|���|���+s���i����q�W�|�W�|-����i���k��0_�U+_��D��F���xs��x��z�k=��9O��W�|��W�|��W�<���7[���+��b�+���__}�D���z��W=��b�N乘�WE}U�W}��W}�;��k!���꣯������ڑ=�P}��qE���L_}�C_���������y>^{����y.��Z�J�������V�j�kc�D�i�Z_{�'�N8�$�W2=��w~�~}��WE=�W���
����W}��W}��W}����S_}��GO���9m>��ݮ��*����
��Z�Z)=������Z)=���N�%s��L_��D^�$1�U>_��U>_��'�N&멯>�꣯�ZO=�Wt�����WX}-��Z�k��Dՙ#Ҿ��Ⱦ�__���n{�?�������J����W�}�#m9Ҥ�ת�k��Uw_{�����^�|-�sd�W~e�qzY��r_)��m_���m_���e�j����
����Z)=�Wt�X<}��WX}m��VJ_a�V_a��G_}��G_}���꣯��y?5I����WE}U�W2}%���竢�*ꫢ�*�k�VO���GX}���ȗ�#����}����諵��G_���,�Z}�W�}��ײ�kY���n{"_�_*m'�n�궯n�궯n�Z<}��W�}��W�}u�W�}u�W�}u�y.����y����W�}���z�<�OC�S_Y�����E}��Z>��2=�GuX������2}��W�}��ז�k��D��%����8��j����Z<}-��������x-�7�_���<��QJ�<���.�<��I)~��W)~���.�+�ȷ��x��&�P&��+:s��WO~����+1�OO�!|�R�O�!�_��'�z�'�z�'�z�<��dz�'�ț�,��_����z"��8��tJ�'�$��^�:�z�'�z�'���k��Փ_=��_��U�_��'��i�HӓO��v�I̯���SNu>�Gujӯ6�j�'��>��CT�~�ྪ�kG�U�O��iB�kG�զ_m�D�U?e
�o9�$�Wb~%�Wb~�Ȟȗw�H̯��J̯��ڤ}%��&�+1�z�'�z�'��+:�,׾��k���_���M�W�~mҞ�C��Q�~��W�~��W�~mҞ�C8��W�>�7�a%j�ȣ:������`�
�kQ��_����_�������'��4�U�_K��6���}m��
�+W�r�+W�r�+W�V�_�����կ\}"^ކ�8�����'�\6|_����_��D�	����_=����Z�}e�y���Z��|������������}�W�}��+����+���s9'd����k����{"�圐���C���
����Z�}5�W>���C����}e�W~�OCJ��J��J���Ӌǯx�Z~���j�+1�V�O乜_��k5��_K���Wu~��B�k�������}U��
�:���k��U�_���M�yz�s���&�+W�r�+W����M�6i_m�����H�\�j����Lב&W�r��M�B����__��|���9/����6J�?�x����> ��s�> �ȣ�Μy�ߙ�"��;M^���&/�~̋|��i�"���紉~�^��Ћ|C���E����E��w�����;M&��&/����y�~��D���^�k�>�ȗ�}Ι�w(�Ȼ�;^��ċ|C�OC�>���s�>���+�1`~��^��!�9��q.D���_��qz���<�3��"_�C=���9�SO��q�E��c��"_�1��~�oۙ��~�Wt2�E�"�N&(�����g���_ ���i 퉜_ �y������mG�/�N8�0�/�m;�>GU�/�=:�>G��/��L/��/���x-J�_��k���7���=��){�o���~�/����g/�N���|yG��/�~�~�z�WtN��_��ik��?��]utP�=��~�"���Y�D��<�c�=�3��"����/�\���^�~?��ȣ:�(�~�G����D>-���E^�G2���8��E���"^���i�q�p~a�_��r�HÀO䰢I�E�?���'���"߶5b�ȗw2�_�!V�_��s��p2��	�"�
gN8s�G���<��o�_�p���'rtP��"߶OC�yE}�/�\Z�_�Q}��������~�À���r�l��c������~?���|�����E^��������Wt��_�}$�>���<�Oi��y�#u�/�����CwO�H���E^��(�����>�l'��E��Gz�_���)�"��H��ȣ:���/�\�/���<��O�"�J[��8R�E\1}آf|"g!5�/�\N9<����[����+��s����9~���E��l�_��,�:�WtRY�"�,���E^��G���|�>��D�/��������o�YH?��<���/��G���|-G�E��Oi��i4����c9��/o�"��#Y��w>��	�"��dB���s9����O�x�y���/��!�����_���qE߶c�2�y��,Z>a�_�{t~a�_��;� �/�~~���E^љC���|�>��
�"_�1���љ�~/O����"�{"}�7�8`��/�9s�3��"߶�9P�y�	e�/�:M��/�>���'�9��"����E�ߒ��_��n�E�G�E��<�H4���s��.(�DN&��_�v2�'r� �_���������_�������C��/���9��O�Bw��s9�h��p��"��-�E��a�~�G�i���yT?��<�"�ꔣf�E�]�O�cT;��)W�G��	��"_�g&l��|��/���|yg,�E��������LԌ��s���/��_���1���ab�"��g>���<��O�"���ŏ)�"��u"�_������M������"�����ț���9Q�/���B���<�O|��yT\�E�g9��'r�Q�"��H����[�S��/��>�A�'��#��E���HI��<����"��,�7�E���W���~91A�/����y����s�Dퟂ�S�
�O��)�?��`�쟂�S�4�O�x�(I��`N��r����ǔ�hD�Wd~}:��F�y.F�'���@~"��H��?���$�i�?Z�_���맙�4�f�������s�!�������;���G��|�L�Ol���?e��������~"��H���-�/�\��Ol���?��'�������������Z�4��������^�'����yG�f��$�E�)'���s9���������v�y���/�����)�?e����d���r�SNl�ш�"���ݧ�������S�O���Y�p}"��/�>I�������9�$��$���4���Z�qzI�'��$��$���b��v���>�Q��"��R�*���y.G�r�i�?-�G-��<�#�Z�yT�hj�Gu�����"�'�Ͻ�Ͻ��Z�y'|.|.|.|.|.|���v���N9-�'ܟ�+��|��O��I�?:�_�O�)���������4�������E�mj�_���?��D�^��	�?��_��}���p���"~����"�y��/��/Z�'rX�����"��
����B��B��B��B�����G7��<�#���U����y.��������������ȣ�]'�N9J�_�!|.|.|n|�
|�
|�
|.|�����K �K �K qW)��g�Eu�\��DՉ�����������B�G������х�υ����y��1���ӵ�ϵ�ϵ�ϵ�ϵ�������υ�υ�υ��R�yEg!��/�iۑF���|Cί��r��s��s��s��s��s��s��s��s��s�࣠�E���;�>�>w>w>�>��_�����Eܜt�c�c�c�c�P��Y�"�s��s��s��s��s��s��s��s��s��s��s��s�`"��,t{�sU���E���n|n|n|4ۿ�C8�҇@
�_����&��&�����G�������������w>
�_��tֿ�C8�\N�\N��s��;7>
�_��Q1��x���E������f�yg!��/��|�0|�0|�+|.'L�{����+L��v������l�"��,t��s����E��'>�>j�_�Q���0L��@��G����>�l�"_ޏ�.:L���xt���E�������G�����#�݇���yG�����8+��_��������ZN&W>:�_��q��s��s�ᣳ�E^�'+>�>�>
�_��;:��/�]���6�y'���V��V��
��
��
�G����3�}�����0�0|�ѿ�C8`�[.:|.:|TϿ�C8s\���[nHL乜L�Q|.ML乜L�Ö{�K��.M|nH|.:|tֿ����݇�E�ϭ������r_�s9�s9�s9a"o���}��������儉<�#�儉|y'��	��/�㊾m��j��;���8�E��)��/�!>>�>�>�>Z�_���a�V��
��
�������������G%��8�+��	�������k�k�/⮺��v�c�c�c�c�c�P�P�P�P�*0��p2Qv�"��rU���E�m������D���<�3ǵ�ϵ����f�y��D��D��D��D��D�\;�\;��C8�\;�\;�\;�\;�\;�\;��1��s9��D�����DX�,��'���r9a���\NX.',��?~���DX�,[�k����&�r�`�v0��_n",K����M��&²�����DXn",��������D�!�&��o�޿\;X�,�����M��&�D����1X��O�!�����&�ra��?��b�-���	���r�r9a���\;Xv�/��k˵�e��ra�v��1X�,
�U�q���g���|�+,����q��jXn5,k��[�s<�°�&��7,��[˭��
�r�a��0���Qq����r��,��[˭���_Q���E���r�a�}�E��V�D�V��+&�Qw���݇���r�a"����rCb�!�ܐXnH,���E���,&�=:W]���s9j���K˯6�����v�ܶXn[,�-&��n[,� a"��@vMc"��#���͍������˝��N�r'c�m�ܶX�Q,�(&��U�&�_��\�X~��r�b�e
˥���rCb�!�ܐXnH,7$��u�� ,� a��u��,w���/-X~i�rb�1��O��݇���r�a��0��p�-�_m�\�X.M,��`�G1G�;��qT�a�m�ܣX�Q,�&�K˥��|�N&�&�K˥��B^�a��rib�4��2��<����C�{���|y'�_��ܐXnH,7$��u��),7$�_��\�X�C,�!���E��V�r�a�e
�/SX~��r�a�e
�݇����;�_m��j��V���[k;�\tX.:,�+����r9a����DX~�r9a��0��mǐ�
�儉<�ƅ��^�r/`"_���7,���ys�����r{`�*0�/�_ �_G��1��+���B�rU`����N 
���U���r/`���_4���/X~9���/-������}K޿��K���r���_Z�%�_����_*���_*���_��O�!����|�>�X��T�ˎ��|y�J"���P�/��D�i��_~�D����D˿��K�?�W��L����_��%�_���<�"*���_*��,I�� �����Kl���Kl���Kl��
�%�_b��8��~)�_!���˯Xb�����o���,���/e�� ��~"߶�KF�d�KF?�W��G3�4�K3��_���|�> �}Kl���KF��
���L��l�
L��q�I�$I��~���=���K��:�%ɟ�C���ҟȣ:�҂%�_*��7,��R�/��`���J��K����yg��"޶�v0��r<�m�%��,��R�/y��{��c�\X.,� �K �o;X.,��`�=��1X~i�r/`���X�,��`������^�r	`��\X.,��`���U���r/`���U���D�����rU`g�q�0�oۑ��_Z���x-��w",��`	��p	���v���˯6��C8s��K޿���,y��K�_Z�\X~��r	`)���)����uK��K��˯#�ȣ:��҂�^�D�����rU`�*���$�_��%�_���|�>�)��_�����<���U���rU`��������&�>��=�\X.L�k����P0��������""޶��u�%��w,� ��)���*�\X��e����/�	`�������K�?�7�'���/�������~�藌~"_���/e�R�/e����헵�K���K���K���������ȣ��$�_����,�~��3_�C�?��!B�����_����B�����"��d
I~H�C�����B�*��<=�C�~�@��/�`"oSn"_������?�����U �����~H��/�~��C�*���B�*��<�7T�!�I�D^������B�����$?,���D���>�����|��C���>����dv��f>4�a���CF2��̇�2��чf>�`��?�Q��:�P���=��{X���}"�SZ��C������=D�!jQ{(�'�\�!�z��'�<�M���)-t�s�{��'��8�t�s�{��C������=��!W�/ �!Wm�D�5��=T��|~_@���o�	 ��Mk�C�v��=T�:�yX�B���?��!D��+����{�C�>��p�i�C�����a/H���P���<,��yX�B���=��!D��s9���!�C��"��4ѓ��|"ߐ3Guz�?$�!1��s�d�:��C�B���"��'C!z��B���=l���ê���?��!�x(�'򯉣�J�P����!�x��Ö�P��-�!+�C)V���a�}��C�Ѐ�e�a�}���f����!0J��>����D��R<��yE��R<��x(�C)J�P��R<��a�|X=������'=y��CO>���Ӝ�<$�a�}Xc�1$D��C������̱�>��!D;�C�ԇ�!W������z>��!W�z�F
�P���=l�Q{��C����<�#�������=t�s�{X=?���i(}��>��a�|H�C�>��pb�Yvև�����|h��f�ȇ��!}�{H�C�:�йO�{tJ�C�r��<��J�
��T~"O��ҹ�=�a�|�3j�PÇm�!��|�C �ȇm��������CF2���>�Y(�}��C3�ч@>�5|H�C�>����\9�4��|X=�ȇ�5|��C��Ň��!D�y���>�Г��<��xX����|�N�xX����}"O�4����<��'��sI�Cbz�>,�=y�����wh�'�~tS�O��J�P��R<���C)6ȇR<,��x�3z�Г�u�!��D���x(�C�𐅇��x(���P��R|"�������ú���O�k9�l}��D�/�x(�C>���Q��,<d�a�{��C���=�ݡ�)wH�C�"�i�H;D�ay{X�R�r��;�ܡ��v�����}�a�{��R��m�M���v��'�>����aS{�����Z�M�!��uȯ����_OĹ�`;�C��찃=D�!�k�C����m�n{";��a�{H�C���=,o��'��/Yx��C���=d�y.G���a�{\��<l}��C8�T�y���!W�z��C�r�ЦO���P�:�yH�Cb󐘇�<��ay{��C<>�Wt���)~�E�V�o+޷}�[<���[<���������-��C01��|��%�[b�%�[O���[)���[)�5�[��[�������޺��޺���v�o)���}����[�=�o�1����-�ނ�����m-�D��)�e����-�6�oY�D���6�/���v�o;�'�=:��`��� V�o��7}ۛ�5�[ݽ��[��u�[~����ZE���|�O��'���o)��ro)��ro[̷��[ݽ��[��-#ߖ�o��ioa�Voa��-|[���۶�-����-����-���;�PdoE��_o��D���a��VdoE�VdoE��_o���Zo����{K���ۆ�-����m��Vo���{���z��'⇦��6|oa�V����|"߶�>��<��Jk���[k���[E�U�[E=��wX��%�ۆ��+6|o���Zo����{���dzK��dz������V�m+���{[����������-��*ꭏ��mo1��9o��9o��9o���4oM��4o����y�O0j�m���I{���y۷�����mo���}�[�m����<�C���-�ޒ�-���譏ޖko˵��zK�'���9!��6iok����[2�%�[2�%�[2�%��&����xے�-�ޒ�|��fO��9��-���i��<��&�i����+zW}��{˯��zK��dzK��dz"O�R��{�yH���[�-��b�|���-s�2�m�V>o[��z~�m�M��[��m��?�g[����[�5�[Ӽ5�[Ӽ5�[Ӽ�[���[������-`������[Ӽ5�[��-��uo�0o��'�m;�����-`�j�V�j�V�j�V�j�m��0o뼷�yk���y���y��'�9����+:�,����i��-`�j�V�j�-M���Cޢ�-:ޢ�-:�r�-'�r�-'޶ro��Vo���o���}���>���}[���۾�-:�r�-'���m���o9�{"ߣ�ľ���fok�'����m���\{[�����vdo;���yۑ=�w���Ȝ��y˜��yۑ����vdo}��Go}�Co1���z�����[N����z�0�r�x��So���]�yE���x+���x+���xˉ�vx��*x���*x���*x[)=�?41���J鉼�@(���[�U�[�U�[�-���-�z߭�ݖEoˢ�*x[=�W�����y�}\�o9�o���vx"�v�lb=�O���9:�m=��&oi��!�']�����-�ۖ�-:ޢ㉼�3G��u���Cj�V�j�V�j�V�j�V���-M�ȣ:��[���[���[���yT����y�E�e�[�m�ޚ�m���xz[<�����魏���-��b�m=���zK�w;1%�y.�c;��q����z��U�[X=�/���_o���Zo���9oK�'���!��9o���4O���2�i�V]o��9o��9o�0o�V+o��VO�p��~��[a�-��bo9�o9�o���x[O���[;���[;�-��r�-'N��Sa�
㴞:E�):N�q*��&U��
NUpJ�Ӗ� ��7��Nk�S�����
O�!
�N�pZ�r�<�#�Nr��St�����8Eǩ0N�q*�Ӗ�T���):N�qZ)�
�T�P8��N��S;��ቼ�̯�e:��i�tʉSN�r��]�iu*��z괞:��Nr�S��6VOĽ��:��Ns
��z괞:e�)sN��z�<�C�z�LO�Q��*�T>O�t�)�S��2�T+���)`N���.�9���i�tZ<�b�C�:��)`���r��S��j�T+�Z9�ʩVN�r��S��:�:�|����!���i��D^�1�iN��S��0�ri���艼�3g9sl�Nk�SӜ�扼"�RӜ��0��9�i�tZ)�2�9��ө|��C��e�D����f��4�e�iY�D��Vb�C�:-�����\>u�E���e:��K����G�>:��i��D�^����G������i�tZ��̱,:%�)�N�sj�SӜ�洧9�iN{�'��	�s*�S����9��9e�y'��&�NˢS����GO��}f
?�Y<�Z��Z��:�֩�N�S~���_��:��i�u*���<�#-|���z"�곜<5�yW���Ԁ�<5�qYx��S���I{"���<5�yE�CZ��J�T��R<��y.��!p�)s;�U�'O=y��SO��r�R<��N+�'�>�m'�}�i�vJ�Sb�󔘧�<%�i�vJ�Sb��m��<-�N�yJ�SO�6i��<��'O=�D�m�T�i�v
�Su���o;-�N!z
�S����8�=-�N!z
�S���#;U�:O;�'�m;�$�)1O�Sb���Kn�vڑ���T���<U�)1�t2��SO�z򉼢����T������Ru�vd��|�?��_ G�6}"�賜��im�D�U���٩:O�yڑ�B���٩:O�y���^딘O�{T���<U���C8�����;a�u*�'��N9Q{*��������)jO��S��f��=E�iGv��S�
�T��\=-�N�SԞ���#;E�)jO�z��'�:s��)DO!�D��cH��B�<��J����Ԧ�6=��MO+��
�o;��N��S�>�7d�vڤ�j����q2��S�j�T�O�r����N5|��S�:�Թ���)}��7�Ӑ��)�O�|
�S ���|�> �>��i�v�4�O�|
�S�������U�)}��4ѹ��=��N�{J�S��������=u�sOk�'������=E�`O{*��&�<�F��m�s��r	��
��̧f>5�y.��@�OF?��pX��>�ȧ@>�)�O�|�����ȧ�=E�)j�'�Ag�\=��)DO��'��I������}�)1O�y*�Ӿ���x<��)OYxZ��Vp�R<e�O�wڷ��o;e�imvj����Ԁ��;�ݩ�NuwZb���|��;��icu�X��O:���ˤOK�'���ԡO�x�2���<���5�y���]�)OYx�����T�O�!
O�x<��O�xI�K�]�GO���%�.�w	�˖�~�v�2=��`N�R��.��D�m�I�=��_���x���%/��D�O'%�.�w	�K�]��Rw�n�t��������%�.)wI�K�]R�,�t�etY]�@�����e3t	�K�]6C����ݥ�.uw�]��|�����et��'�Y)]�3G�]"�R�t��9`D�%�.�vɯK~]���Z�ֺ��%�.�'�<��%�e�uYb=�w����m��d��z"_�'�����%�.�w	�K�]��|����9�4�e�u�X]�S����ݥ۞ȗ�NI�K�]R�r�-�e�tI��J���!�.�v�K�]��x�D�%�.��D�/Ev)�K�]vQ�]ԥ�.��K�]"�x�D�%�.��'���v��K�]"�iO�V�����y.G���.xi��^뒅���%�.�w	�K�]�9>��B��	��eGv	�K�=���)�/xi�ˎ�Ҁ��4�e!�D��hmv)�K)>��p<��˾�o���e��D�����}ۥ:/�y��'��|B���ļ�۞Ȼ�HS������'/=y��K^�𒅗��%�.uw��K�]��Rd�"{"��Rd���������SɯK~]Vp����֥�.uI��r�RQ�}�e�v	�'�
�KX]�겕��֥�.�u	�KX]�겻��֥����>���]Z��Z���ew�D��|pSd�"�٥�.E�D�	�exI�K�]R�r�H�,�.Ev)�K�]��|C>l��]��Rd�"{"����H�_��z"ߐ[���"�٥�.��K�]"�i�H�l/�v�˶�Rd�"����+:m�.Ev��]��_����֥�.�ˆ�_W��Rk]Z����y?e*�K�]���ZO����.a�D���I~]��_���,�.K�'�\>��#M�]����tۥ�.�vY >�i���m�n�tۥȞ��i�m��.�v�K�]��_�ֺT�e5x	�KX]��-|"ߐ�|��Z���%�.�uɯK~]���%��ȟ�OV��i�H�D�%Ҟ�s��eyI�K�]����{"�蔳�|��K�]v���{"���m�n�tۥ�.�v�'�F��f��D��)'�����x�/��D�81��F�8�x���/�x)�K)^6��,�,I/K�˒�|�~b��x|"���<NL��'�\Q�y��Ku>���ϵ�Q�:/�yI�Kb^ֲO����Sb^�ғO�r<g�ļ�`/;�'��G�K�^B�����`/�z��Ku^��R���,\��+:���%1/���F�8�ļ$�%1/K�Kb^��9��KO>��pXI�Kb>�W��8�$�%/�xY�^z�ғ�����'/=y��KO^z�ғ���e�zٮ^��R����eozi�K�>�o�a%W/�zi�'�=�x�`/�zY�^�����%j/Q{������7��M/5|I�K�^����O�|��J}D9���lW�����'��b������e-{��^����$�$��q.o������<��������ys|.�����s���@�*P�
��e|Y_n���stl�PP6ȗ;�A�=P�ʗy'�;y?o[P_ԗ��rB��Pn"��y�1-�/7�M����\;(����r��D(7���c���cg����XP�j8n5��[���r�D��z�W8��W�+��c��q�a"��\=��O��C���3}��z����qC�!q\�8�C��]��.�c��D�=�VL�!���Պ��q��Gql�?�V�(&�����ܣ8V�O�!��m���q��Zq\�8�V���Պ�j��Ǩ��s1j����Ʊ^�X���8.`��'�'d��q��ؒ\�����/�;�����qM㸦q\�8�w2���yg��ǖ����q�mq,�?.`0�]�ǝ�c���|��77����yz<.s�9���e��2�qs㸓q��8�d{�����͍��qMc"�����2�qs㸦q\�8�i��kqW�埈[�2Ǳ����q\�8v�77��qW��8��4�kǝ��Ʊ8���q,�?�d��kǝ�cq�q㸀qܶ8�QL�-t��Gqܣ8.M��pi�!qܐ8��[����:ı���!qܐ8nH7$����J���q��4q\�8��c�{�=���"�<�VW+���Պc��D����q�X�\�8.`L�|.`���;���Ʊ����1��p<��q\Ә��k�5��<��͍��w2�_p�r����qs㸹q��8nnL���w�9���/8~�q���q\�8�|;��+Ǖ��2�q��X���?V����[ �-��ȱ���r�9n��@���y'��.�C����]�c/�����Qr,�?n��G��#�����q1�r\9.�C���Ǖ��~�q��إ���+:-�?���@�[ �����q���1�/�,t���q\�ȷ�3���^��2�qs㸓1�Й�0���-���Պ�e�F�	��{�=���q��4q\�8nH7$����f���q���Y�?nH7$����{��|��t(�Gq��?�VW+�{ǂ����J#��GK友�R�גn�����u���ñT���p\t8.:���6�c��C5�N�1�݇���+V4����ǭ�WVg��9�C�!���݇��q���p��?6�䏋�E���q���p,�?.:�[oy��C8s�}x;�F�'�m����ı���oy.��K�u��V�q���p�jx�5F�{�M\txB�ȑ��q���p�j8n5���
���r�q�cp\(8.K�;ǅ��B��z��*p��M��O:n��2�N&���ǽ�c��q	��������u�G�l�?6�-���䏖�=���N -����⏖��#�(�����A�h����G�T�yE�M,���+�[k-���������T�h�'��;`���&�\V�����U���qU�*p,�?������%���q	��3�?�
K句�G����7�HS���Q�y���-���-�D^ё��?������!���I���I��T���J���J"��K�T�G�T�ǂ���?*��<��K�$�G�$�G�$�G�?���<��K��GY��GFd�GFd�GF,�?2�#�?����?:��s?V���ѹ��ѹ��ѹ��ѹ���K�إD��J��|�N9Q����8��Տ\��Տ]�G�~�ҟ�[�Hӹ���^�Hߏ����'��/Q��q��`o�z��[��r����m�o�z��[��r����\���-Wo�zk�[���8"O�dj�x��[)�J�V����-o�x���^����%�yz��Zu������-Do!z�[u���R|"O��jYx���z�Vw����ܭ۞ȗg��]���nuw�����|��{"N/�n{�����|��{"ߣcH�݂�|���ݭ�n�v����r�%�m	����|��{"�dRw��{"o�cH����Vw�����o�v[�ߺ�Vd�"{"����m��RK�'�< �����-���a��n�v+�[~����qX�?�k�q��ן�C8sD�m�~���z��mO��&�����VK��.�Vw�����-�n��[��R�rO�v�,����-�n�v�l��ط"�٭�nk�[��"�ƾEڭ�nEv+�[�݊��	񩩵�mg}�F���L�d�%�-�n�tK�[2ݒ��G�>���-�n1t��'�F�Yߒ��G���-�n}t+����CO��;M�ϭ|nk�����G����-�n1t��'�:���o�s�cH��2��4�Z�����!;�[�ܚ�V+�4���mA}K�[a�VϷ��Cnr��[tܢ���q�q�����!��9���ƾ��m�}��[��:䶠�-�o�[��Է4�m�oir���6��!��u�m�|� �
�Ͻ%����'��D�mj������|ێ����톟ȷ����Vn��'���[����d�|� �6ȷ��Э|n�s+���V>�u�|n�s+����A���y.'���Uԭ���sZ:��֭�nau[P���N��>z"߶�ʞ��g�-�oK�[X��̷ֺӑf�|�3ߊ�Vd�����-�n{��R��T���yE'�ֺ�֭�n�u�[X���V���y'����_����n{�[�݊�<��Q��"�i����۞��J����r���ˉY>�	�'�\�G�w[*�Z��Z�ֺ�֭�n�uk�[k�����-�n�[�݊�Vd��mA}+�[�݊�_w�1Pk�6ȷ�-�n�[X=��1��n���Vd�"���m7|[������nEv+����i�H�m}o�v���R�r�����-�n)wK�[��R�.���o��D��G2�'���&oK��R����ļ%�y.'����-Do!z�[�ު�V��u��Z��Kb�󖘷�:����xT���:��+�,g�|� �6ȷ6���-Do��D^щ)Do!z��[u�z�֓�x���m�|��'�mK�[O޶ѷļ%�-1o�yK�ۂ����U�:o�ۂ�֦�6���:o��6�֦�6}"��ƾE�-joQ{���f�����y.�ϵ
����m��ȗw<��P�>���QQ��:����-�o�{��[��:�n�1E�`o{+�[���̷��E�-joQ{��[�ޢ�����E�-Wo�zK�ۦ�֓��|"޶ļ��'o=y���v��J�%�-1o��[b��V��,�e�m��D�]���]�m�y+�[)���,�-6o��[<�����PP��R�5��ȷ휐��,�mDo�x+�[)�6��x|���_��U�_Y�Հ_[�g�xE}�,��¯,�j����Z ~-���k5��|"��P�R�+�R�+徺�۾��+Ҿ"�Ȟ�C0`�'|C��Z�}-�u_���__��'�~1�"���}E�ע�۾��۾Vp_)��r_E�Ud_���Z_��'�ʯ���E�W�}�W�}�W�}�W�}��r�k��i_��i_��i_E�D�	�M���W�}�Wk=�o��a����������������~}U�WE=�Wtt|<O\a�VO��;',ľ*�|�<)L�vNh�'���*���W�}-ľ"�+Ҿ"�8�n�궯���r�۾"�+Ҟ�+:s,׾"�k��D�ɤ۾��Ⱦ�k_��|&�=:`t�׾�۞�s�&�\+��������+��y_��U�_�����Z�=�����D-����_��Փ_{����Wb~%�W<~���y_��D�/�����=��r��~��6|_����_����_����_��'�\���_!��_������ί����}U��
�+D�B�+D��r_m�զO�p���o��&W�r��:����x���
ѯ�W�~���V�k+�U�_�U�_��'�\�G��չ_��չ_������ܯ�����>c��}�W ���s��iw���O���@���j�k���_���_5�U�_5�U�_5���_���_˵���*د��Z�}�ྡྷ�+j�
��`�
��V��������_����Z�}�yT�۾�m_�����n������~"���v�)믌����WY��Jl5�W-����s����`�vw_�U�_�U�_�U�O�0���M�B�+D�B�k���_��6�Z�}��kw�D�B�l��
��`���_Q��_��_�¯6���=�o�9a���_!��_!��_{��6�jӯ6�jӯ=�Wu~U�W<~����������+����+����+���y_u�UwO�!|\)?�Y�}5��C+K���~_K����y}����k5���_����_��զ_m��_��U�_��U�_����
ѯ�|"��Ӧ_m��-��կm�y.�������`��O��r�H��_!�D���Y�կ\��կ\��)~�ך�+j���+j�
��M���+D����:���:��+:���W�~U�Wu~U�Wu~%�Wb~��W<>��p�I̯�|"�#Mb~%�WO~m1��񉼢cH)~e�W~��2�k���_Y�=��U�_+˯x��ǯx�*ůR�*ů��W<~��W~�'�J�k����Z3~5�W�}��N�+��R�۾��۾��+Ҿ"�+Ҿ������__���__��D»��Pd_E��S�j���׶�k[��__���-�*��"�*��"�*�'�F;�,#���_��i_E���������ʯ����N�Ⱦ��ȾZ뫢�ȗ���}�V_a����~U�qE{���c����ɶ�k��m_��'�+u�Uw_u��@�
�'��~��_Y���O�iב&���k���@��¯�W)~��׶��|�N9=�Փ_��D��i��/��U�_��U�_��U�_kƯx�Z ~e�W~e�W~e�W>�w��(��U�O�s�W)��Q#_�w~��+��m#_�wX�ȗ�V/���Ei��V/�D���E����E��wX��s��y�ߏn/�~�>���s�~�{����r���C���y�ߑ�"�����"_�wX����;�^���;����
�=��'�y��G�y�������ѿ��z�w����E�w<��s��ǉ~ߋ<��H{�/�ȿ�+RY�"�oF�"��,�ѿ�C8��/��O|9D��/�\����9�?_!�!���y'�`�y.'&�~"G���0|CN9Z�_�r�Ql�"���܋|C���Y����rb��W�x'|X����&r��u�"�������ğ��
��"_�a����߿�C@�_�ۆ俈C �_��;���/�mS��"߶3�F���/�G-�/�N8 ��{e|y�@�9��/�
���qEO����E^��p�y��C�_�k��n�E�!��SY�"ߣCb�"����	u>��O�"�s��/�\N z�����D�����c�_�Q�R_��Q�L����s����E�U��_�QV����C�4W��Ʉ:�����Ӌ�_~�C���C��M�o��GI��<��>��yW�����dD��r<b�_��W��O���yg!��E�!g!��/�=:���/���[�C���;D7��"NOS��8=6�}E�G�3�v~Ѯ�"����/�N8���/�=:Ҁ�/�:� �/��zsVx��-{^�ɴ�Lx�y���E��[���C8� �/�N&Z�_�_&�6�E���B��<���p�yT����n�yq�/�>R�"�xȿ�z�mS��"�Wȿ�C8���/�>˥����y.�#��E�/�#�/�\���+��E���`���������Y�"��C ��/�Z����9�U��_�|D��+:W��/�Q�����B������0��tÿoh���aE���8��E\Y�"^���yEg��E�1�����#��E�1T�d�����ߎ���[2�����nh���C �y.'f�E���B���<����y.������Wt2�_�!|T��E��ˑ��߫�Q}.Dֿ�+�,G����f_��E���<��w���|����C81!�/��UH��8*$�E�R�q.���8�/�F���<����"��\�ȷ�\��E�	?�_��X�yT2��EէG��Ddx��<�����Yݗ���ǹz|.<�ZJ�_��Q˪��<�C�U��|����ȟ��w�����:����O�����;���/�㊼!x��8��E�?Z��_���)��"�dB�O�b	�E����>���>���"ߐn����T���+�HFo�D~�k?��_��k��� (�y� ��y.��P����N���<���"_ާ!H��������"� ��E\3?��h�q���ܯ�ܯ�ܩ?���N �_�Q����G�A3�"���̿ȣ� ���Gu��_��C`�yzW(o���!��E�!gf�E�/��ut\?��'�C@�E�!�u���>��&t���+�9���y�C��y�s��/�=��s}���_~%��c�}����������������4��ȗg�}��Ol���?��'�����?&�'��d��f����E��0�����T�O��O���?5�G���<�i"�#�����O ���?���s�D��?̧`���6�Ӧ����;�����}�/��0M>��`��\�����O��}<Y}r�O�>�Q�����"�j�?���'��e�w���O�}N��牏�y'
z�O<���?����4������.�d�,�����O�P���E�<�7����/�N���'�m;`h}���Sӧ:�T��|"���ѦB�O��Q��"^�>��Z��D�!��G���<�3�>�qWU�yE�M�s���[�\����E�`���\}"_�aE��|y'��/���=��i9���U�/��}6Y�!�GI��<��I��i�?�_��;h1�Gu��?���4��|"�(�4����|O�
��O���b�"_�O'��O��QF�"ߣ����J�2��%�'�4���Ӏ��O��	�?��D�G焺��S�E^�')�'���ܟ���r"폶���>�H�?)�'��(�~�/�S=�/���!��ߟ��Sw��O��i�?�_�ttl?�h�?�'����M����ql��/�9'�sb��J�'rN(�?J�_�!�&"����&"�O��)�?E����ٟ"{>�y.g�H�i"�OX��?1�Gw�D�M�i�4�E�/�m;��~�W�sG��M�'`�(�~�0�O�����"��4��O����"O�C����92�O�<�WtX�O0����������4����谢�E��ɤi��+:�4�yEg�Zy"_���'`�̟��0�O����"�H�@�E����)�"��5�/�G딣y�E^��'�������$ӟd��L��O���?j�_ďV���?��D��$����y��Cb�O���"~�b�O�)�?��V��ʟZ����E�/ǐ4��&��O��I�?i�G������/��WN�r2��I����?��'M��ɟ4��&t�O��!��ON�i�?��D�^;<G
B�O<�/�̡��E^љ�
�T���� ��O��)y?%�����E���#��d�E�/�!%�����~��v��O������?^޿�>�P��"ߣ�:�y��94|�����
�ȣ:�(�~������1�j�y���Jt���?��':�ڑ&:���y�E\��_:�O���?�C�tȟ��!:�<��Q:�O���O�"��xT+4���s��%`��C�������>�O�"��/��П�Cb�O��ɜ?��i�4͟���y�E�	'����4O��T�O�x���E^�Y(s���S���yz?^���/�ԌO��@1�'���П�Cb菚���9��O����?i�����C�>3]����~���r�V���0��}�/�>3��?��':�Dǟ��StwO䣏v����E�!�!�?U�
�$��xI�����b	�'�=�
/��'�\�%^Bቼ"`	��*x���x�����^Vp/+���xi��vxٷ��񈱴�˾�e��R/9�\{ɉ��xɉ�M�yE�вo{ɉ��xɉ���yE�RO�{�c"��'�e��D��G��V^�m/i�6{"���Zj�V^6i/��!/��!/�D���&/i�{Y��t�K����^��%M^��em�R+O��;�,�^�e����zi����0/��R+/��D�!}��y"��d�#{Y��,�^b�|^��%s^���xy�H�B�e��R>/���4���eG��4O��L�%`^�%`^j�V^6i/�0/���M����|��s)���y	���y	���yY���K�<����KӼ4�K���K������C�+�����g)�'�\|���s9��Т�|^2�eQ�R>/��{�ݽ��K=�w�a%�^b�%�^b艼>YY��,�^�~/a�V/{�������e��Rd/E�Rd/E���{����ˆ�e��Rw/u�Rw/)���{I��u�Kݽ��ˢ�%�^u/u�Rw/u�Rw/u�D^��(�^���q��g��|�����K�=�Wt�	���{I��u�Kݽ��^u/��|/��|O�|p���Y(�^��eQ�Rw/)��o{����{���H{���H{�ʽt��V�e+�Rw/˵'��'+k���{"ސ�{Y��,�^6i/Y��I{i��|i��|ٷ�d����&��eQ�R�/Y���/����{i��|i��|����{����{�ʽ�K���V�e+���{�ʽ��^6i/���I{�ɗ�|٤=�7Ǒ&D�ȣ:���K��T�Ku�$�Kb���^��:_6i/��R�/����/Y�|/u�RwO��5|�4�����R�/��R�/��R�/��R�/ۯ�,|i��U�K�d�K�d�˪�_�_/ۯ�x|Yu���y.G��|"��H��/����/��D��'_�_O��;����'��+�[2��D��g9��R�/��D�7!��/뼗6}"�Z�G�D�^���ˆ�e��/!��O�����<�CT����K����yW�B�e���\{"߶㱜rB�%D_6i/���\}�՗}�Η�|�Η�|�Η�ˎ���:�l�^
��`_
�U~�\{)ؗ6}i�'���/ǣ��K��l�����/���z)ؗ�})��q�(ؗ�}Yb��cH����K���^��e���/!��Rzi�'����D�G?R*ؗ�}YO�D�yT��t����%}�ȣ:��K ��^��g����/���/�R�/5�R�/����/��D�mG�~I�'�\N95�R�/5�R�/+��@~	�@~	�@~	�@~�ʽ�K ��K ?��/���@~Iߗ�}Iߗ�}"�곜�}Iߗ�}Iߗ�}Iߗ��yT�~��~Y�=��r�
��})ؗ�})ؗuޫi��t�K�>�/����͢�`_���M_����/��'�=:���^vw/Q��/�D�h�9:��s_V�OĹ��q'�K �l_��/��R�/5��/��'�9��e��R�/5���{YԽ,�^�r/��D��[2˵'�>F�藭�KF�d���̤�_2�%�_2�%�_�%�_�%���C�e+���{�ʽ��˾�%���?��}\�\{)뗲>��!�˵CF2��чܡ�e�D��+����C����<*�)$�y>e�p?��!��~�C����=��ȣ2������?��!��s�!6���[Ȩk�ý�p/ ,��N�p/ ��&����4����6���Å�p� \(
�p� ���Å�p� \(��F�p� \;����p!�D7����$=�W�&⨮0�+�
C��0�r_!�R���M�p!�Dw&����p9!\N�&�9��e��Z�p�!�`���p�!�j���p9!�`���p9!lj��!j�z����k�BAX���;aoz�P���;aoz�c��;aIz�v��;�|�t{ ��&���������aoz�c0��p�,~q.L��֟����@�un����@�=n���΅�p� lWw��p� lW
��|�Nw��p� ����큰]=\(�½�P���?��yzg��?�3G����|�>�,ǐ{�^@(�C���P��������%�����"��?��!�y�D�ϵ.L�|�rU \W�U�pU \W�"�pU`"��sU \���U���~b?��P6ȇ��A�c����y�|�r!������'f81];�&�N�,���D^�g9�&��U��}���>�����p9!\N���x��+LĹ,��b�xgg}���>�[�BXc�0�5��
�D\�{�C���0�5�a�}��n5��
�B���؇5��VC��0�W�?n�+a�}Xc.:̈�/����p�!\aW��p�!\aW��p�!�1w���<�c����|yg����BA�P.�a��D���õ�p� �1�����p!�����p9!\N�'�\�w��p{ �
���p� �1w��p�`"��q� \(
�p� �1w��p� �1w��p� �1�ȣ:�\;w�����~"��dJ��1w��p� �1w��p� �1
�p� \(
½���~"��S;����pU \���6�pU \W�U���>��½��<��]��;��+��\(��s9����J��<��2�!�
C���0�+�B�v����@�.�5��^@�.�K ��;�C���O���TN&W�U�pU 쿟�s�PV���p� �1����Hs� lɟ�C8�\N��儰8"���s_!��W�z��^?\aW��p�!\N���p9!\N7�8�\(
��pU`"�>���\W�.�p{ ���.�p/ ��B�Z��|yG��?��!�-h�C�Z�����!�y��'�\�߇�?����[��%��%?�� &�=:�����-�C�*�P��>,��}��C���<�sBlb�ۇ�>��e}XvÇ��!��}(�CY�Ňu��}�&���T>$�!ɟ�s9MT���I~H�C�����$"�e�}�l?�Gu���������e�a�}�0�Wt	�C�6ۇ�?����+�C�?���9�:���I�Z���?��a%~h�C�����>�-�C������I~��C�-�ߢ��`�r��:ߪ����E��-1��~��V�o����o����o=��~�ɷu�[b�%�[b�%��n���J��J���;�?�m����oY��.~�·,|���{����{K��H{���H{��'�����"�-��"��ފ쭵�Z뭵��ꭢ޶�o��~"���̱~����v�o���_o��Vo}�V>o�ܷ}�[����>���"�y�b�m����}[�%�[2��s�*ꭢޒ魏�V�o�ܷ�����-����ȧ�m���Zokٷ�z����z���z"��c��[�mW߶�o}�D\Q���[�������Z����ֲokٷ�z��'�|0�6�O��r�����[X�U�[2�%�[2�%�[2���yE��y˜�r((���y˜�%�yE��]��b�iޚ�m���9O�_�-�[Ӽ5�[�������me�0o��Vo;ŷ�x"N�C����C�6�oi��!o��o9�o9��O���.��oU�VoķPx+y�m�[ɻ�[}�����o����n����n���lw�v'��;'��8;��rt(y��w�v'�\�Na"����[��e�[��5�[}�շ[}��sBj����N�m���@|[ ��[���[j�����-��R�m[���n���n�·�v"��Q�n��@|��շ[}�շ۶�-��V�o]���n��n���ڎ����|[>�ޟ��ɶ�m[�V�n%�V�n���lw"����n�·m�[ܻŽ[ܻŽ[ܻŽ������I<��p~�{��w�{��w�{��w"�2�m��f|"���So�Ƿ��[<��p�I��xK��x�)���[�Ž[ɻe�[���[���[};�W�1J}�շ���m����n����n����n]�{�j��v�j���
�m���n���n��{"�}9��O`�yo�{"��Q�n��{�j��v�h�bv�c�<v�c��u�W�2u�5�g��Ǝ�m!��n{�����Z�۶xz�2��[`:���h��&���-���m=�V�n5�V�n5�V�n5�V�nQ�<u�Z>�D�%�yE���j�-���m��V�n��։n��<l{E?�HG�ttKG�ttKG�tt�k��ޖXo�鶋zL�]�[s:���#0��C��!Cݚӭ&�j҉<���Lo[��ukN��tL�e�['��[���6� �
�-��BΉ��3��&�Ή|-��[�9�o��v+o!�rn!�D�����yE�!�B��['�u�['��i���-�ȣ�!C`:��wNX�e�[��e����L��ԉ<��pѯn���~u�W�~u+S'�> 	L��t�I�Nt�D'���-���-���-�ȣ��E'�m����}}f��n��D�g&��xzkN�-����d��V�ne�V����Ԝn��D�މi����n���]��.�-V��ԭLݶLO�!��Lo���n�궋z�W�]�[�:�W��I�m����-|��+�߭��������?�%���m����:-�����i�uZb��X���)�M�S�vQ�]�)��C0�R�zߴR:����M�o�}S��G�l7e�)�M��S���� 7�i�sjtS��ݴ�95���M����洧9-RN�mJm�>�Tߦ�6��)�M]m�t��ڴ�8�Nm�h�*�Ѧb6���Myl~<�Lĝ��8���M��F��զ�6m�ț�?d{�S}�R�Ѧb6�)�Myl�����i1p�WS�:�/�ǚ�>8�N�S�:���_�v"��3@�cӮ��¦6�
��C�cS���b6�i}p*fS1������5��)|M�k
_S�:���V�U�iq�hSD���b6�Nm�hSD�"�Ѧ�é�M{�Sj;��rX-�:4�i;q�vS�����N��v��N��O:)�Mۉ'��ojRܛJ�T�7����M;�������Ʃ�M;����8��)N�'��%��Ľi�p�}S�zߴw8��)�M%o*y�b���-�)�M��S�;��p2��B�
�P8��)N��F�+8��M+�2���vx"�ꓕ�8��)'N9qʉSN�� �-�):N�q��St�მ�8E�):N�qZ�����)MN�'�\�4�r��Ӓ�>8��)M����=��� �Z9��iWp
�S��j�T+Oč�>85ͩiN�S�<��rb*�Ӓ�T>��9�ϩ|N�s*����T>���)�N1�D�B�,,NuZE�V�>:��)�NK�S�b�C�:��y'��éiNMsj�'��|�N9ۉS�2�<�nv�:��)sN�sʜS朚�L�,`��+:�5Nk�S����0�Zy"���J'�49��)MNۉS��:��!O��q��sB��V�U�)MNirZE�j崊8��i�pJ�S����|�N�rZ�扼��sJ����>8-N�D^�g&�rZ����&�4y~ؾ����!�-�i�oʉ��ߔ���i�o��St���<���b��&����VN+'��MsZӛ�9����圐9��y"O��C�e�i�o�'�N8`��M�}SE�*���:sʇ�uZ�����Z��:��i�oʯS~���V��:Uԩ�N�D�'����:�֩�N�uj�Sk�Z��Z�e�)�N�uʯS~�6��5��������+�{S~����ZO���i�8�l�ȗ�	F2�v�>:�ѩ�N�vӶ݉|y�m�)�N�tJ�S2��鴹7U�iso
�SX�6��5���NxS~���x���_�=�qz�uS~���Z7�����D�G�n;m۝ȗw�H�SʝR���|��;ߩ�Nuw��S�=���iH�����m�n;E�)�N��D�ɤ�N�uj�Sk���:��ip��Z�8m��C8�lN�v���������NEv*�S����Td�";٩�N�|S��"�i�����N�v��S����<��Q��+8٩�NEv�<�7�Yh�D���PʝR�r�H;E�)�N�S��"�i�H;�N{�Sʝ���m�n;E�y'�U�y.'��;���Z>�I�S�����m�n;u۩�N�v�S�]���mO�{�����ݥ�.u�D��/ۜK�]��<s��|.�w	��艼_�ղ�d�et)�K)^�����ղ���.�x)�K>�Wd�N�!�e�s��K<^�񉼫�ƭ��'/=y��'�Ѳ�,x.=�D�!�\Y]B����ϥ:/�y�����e�si�K�>�7��Y�E���,�.ˢK�>G�R��/+�K _����]i�K3_���?�4�yE�'�|�.e�D�	g��,��$�$���/{�Kl_b��׺��yE�%��9-�.I~I����<����|��B�K�_6V�����/y�D�!ǣUץ�/�~}N9-i�˪���J�T������p"n�J�T�e�uYb=�W�)M�_���p"����������%�/�~�~]�_�����%�/-i�K�_Z���"�唓������O�?�Wt�Y�]���p��ۮ�H�򗖿��yE>����%�唓������%�/-	�����򗖿��%�/��:���O�!��p<*�����(�ʽ�r/�\(� &�m;]({��%��|�>�ʽ�r/��(�ʽ�r/��(�ʽ�r	�\�ȣ:�\��C�xgy�cP���;�A�cP��;�A�b^�
����/;�K�_���|y��⿴���/;�˶�-|"^k;��n*���$�$�%�/I~I�K_��$���y.g�������/e}�)^����O��9���@�����/}	�K _��f��/k�KF_�i����C8`��%�/�}��Kl_v��������/�����f�$�%�/I~Y3^֌�p���%ܯ�#���,#/I~���2�䗲�l/��'��}��O�-�їm�e[x)�KY_V�O�{��ʶ��<�SN�_*�R��N��1J�?���1J�_�������e�x�P.�K e?y�P.�K �@YY^��W��Q�_����������C��R�_���<�����r/��([�˽�r/�,6/[����xy[��U�rU�\(W�%��f�\(;�K�_Z��򗖿����/��'�������/�~	����|-����?��{tN�P��R������e�yi�'�N8M��e��D��!�/��D�G�rtخ>�7���@�P.�����/���K�_������"_�ѡ�/�}i�K3_��O��k��
2��ї���%�/�|�O^���̗e�%�/��KY?���y��䗕�y��J�$�ee�D�/�qt��K�_*�R�J�T��ҟ�s9:$�%�/��K�?�W�c��l���D�-Y�^Z���U�3�=���\(�)�'��4� �%�����(�J�?��pZ�^��R���"�H�2�ʽ�r/��x/� &�NL�ʽ�r/�,�/���U�rU�\(�ʽ����,o/����r{�\(W�U�rU�\(W��r{�\(k���r/��(����r/��(��>�rU�\(W�U�R�O�{t	����/�Y�^���p���e�z�����R������/y���:��e/� �%�r	�\(�)�K�?�WtX��K�_�����������/-i�K�_Z���p�T�e-�D�m���%�/y��˦�R������/y��K�_��#�?��#�?Z�#�?��#�?��-���������G��s?Z���?Z�c��D^��y��G�T�G��Glj?b���?6�e�D�����?6�������D��)w��G���>��<���'�\��_��#�?��c����-�����Q�e�Q�e�D�Ue���K双��菌�����d����g�������(؏�G�~��?
��`?
��`?
�#W?r�#W?r�#D?B���4�/�Ц��m�y.��\�hӏm�����M�Ȼ�����'���]�~��?
��`?V�Q�Y>�(؏��G�>W�z��ڏ��(؏=�G�~��G�~��G�~��Gu~,�?��m�Ѧm��!��!��!�����A�я��������:?6���Gu>�WtX-����y����Q���Q�{����Ώ���ɏ��G)~���>��?J�#?��c�Q���р�р�р��'�m+�O��?v����h���h�'��#�>���>��#�>��"�(��"���~�yz�D8'�G�}�Ǌ�c���m�܏}��>�cy�Qd׏��G�}5��c���r׏�����#�>V����mOďc;:��G�}�R?R�#�>R�۞�C�c��Qwu��J�����X�~��*���>���>6��Ϗ��G�}��G�}���F�#��s9���G�}�R?��<��+ۏ[��c���J�����qE�}t�G�}t�G�}�G�},I?����i���7���>"�co��7�趏n�趏U�G�}�R?R�co��7��'�\~t�]}"�SN�}��G�}��y�����������~�����?��>R�#�>���>���>��c-���}"���Z�#�>R��>��|y'�����~T�G2}�R?*�c��V�Տ�����%���9��>�PQ�ԏ��؛~�M?Z룵>Z�#�>��#�>*�cI�Va�D��O0�룵>Z룵>Z�#�>��c��)�mk�'�\>�(����ȯ���خ~��*�#�>��c���_���_���_���ZO������#����-���+*���G�}D�G�}��v�c��D^ч�ԏU����#�>R�c���r��i������u~��ys|��r��dRw���m���_O�r�(��"�X�~��G~}���*�c��D�˙��>Ǚ#�>R�#�>��c��i�ԏn�趏U�G�}��G�}t�G�}�`?���>v�)�i����}"_��$�>Z�#�>��c���p�ȯ�/�wՑ�>Y�����G�=���N8u������>"�#�>���ۏn�趏n�趏n�(��}��Z��|-ǣ������H�'��8�$�G2}$������>*�h^�1$�>���xy��u2	���������3|}-ǐ��H��>�裏>�裏�����#���C8���G}�����>���+�̑L��D��SQ��4�N}���H��d�H��d�H������>Y)����(��-�G}l1��	������������������������������[����ؼm1o1t+�[����V>��-6o1t��ۮ�V>���|n[�[����W��k"�,l[���VQO�O�)�������h���V������-sn��D�{��Z���V+�Z���yE�U�<>�7��՚�<OV-sn�s[Y�V�����mey[Y������Uԭ�nk�[2ݒ�C���Э|�ȣ���v����q%�mx�������%���|t���!�n}�D��-���C8s>g�ֺ��yT�Z~���<�ZX�*�|y~��V������m�w����V�����-���C�0��_�����-�n���_��m�x��[��������m��D^�a%�n�v�)޺��m���m[x�[�݊�Vd�m����m>���Uԭ���?����V�L�E�-�n��[E�*�VQ���m�n�[E��y���U�mww��'�+au[���yO乜_����-�n��D��$�v�#M�=�e+�D�A?�)�[k�Z붂���m+�D^�O`�rO乜9��λ��-����dRw�����n)w�����Vw���m+w�[u�E�-oYx��[>�Gu<��[<��񖅷,��ϏJ񖅷uޭo�x+�[)����=�mx�ޖ~��U�'��C��&1o�yK�[b�֌�꼭���n����-W��\���Momzk������U�'o��[)�J�-�m�������'o��[<������mx��'�=:s4�m�w�������n�����ր���-�n�vo���ڭ�nEvۤ�6i�n�E�-Ҟ��ewK�[��R��m�n�m�n�v��[�ݶr�H�E�mww�[��6i�ֺ���}��Z�����m�v[����\�٭�nEv+�[���f�H�E�mm�D^љ�۞�C��(uw���
�o���y}�-�n˵�r�\�-�~_~n�!�rVp�����'o=��Jf#N_Q��:ﶻ���n����91ˉ�`_�h�!|f��u�so����y'����o5|�����ȿoA2��m��[Fߚ��1F�˱]�m���#��ض��%���o�}��[����������F�I��oe}[l�b�ۿf`"(���Z��C8���-�o��[���������o��[����߿v4#���oK�[����߷��U�y��q�Z��Z��Sb乜�����`�p<�������m��;���mS{��[���������-�oy��ފ��򷖿��m�z��[�������-6o}��[3��ȷ��-�o�|��b�ȷ���m�y�O�j������l����] ��������mo5|���2���f#�����u�m?yK�[��V�����-}o[�[�:����-#o�{[F�6������my�<�����7䣏f�mo}��[Fߖ��������oe}+�[Y���O��\+���C8�����o�}��[���$�-6o��[�����|-�$n�����o��D�5�뼵�-�o�~�[����������o-�[�ߒ���|"_�Y(�o�~��'�=�1P��*��żm1��+��Z���$��,o+�[��*���|"ߣ�K�ߒ����~"��H���������<~��W-#�������������F_;ů�WY��W3-��+��ve�WF?�o�1te�WF�'���k�D^�G�+��2�k����ZF~-#���+ɿ֌_���f�����������'�􌡫����+j�
��`��~_K���}"��s�:��s�V�_��չO�!��w��yG��~N Q��x�:�+j�ȗ�߶��Z~���j�+}���+}�:�+W�r��|y�m�>��O`W�~����+j���k��D�G'�ǳ�U�O�k�<q�W�~���,��r�k[��-|"�ѹ_��չ_Q��_Q��_Q��y��<~m�j����:��s���_��չ_Q��_�ɯ���گ��W�~����_��-��~������G����#��_��U�_5���_Q����Q�O�k� b�U�_��D^�a�`�r�+W�r�+W�r�+W��s9�����k��O�Q��W�~���j�+D��~_m�զ_m�զ_��Փ_���_��U�_�ՀO�k��]~5�W~����+���+����+����+����+���+:M4�׶�+����u�Uw_)��m_���|"_����__���__��Dܯ��>u���H�����yE�n����m���}���~�F�}��V�_�����
����
���yE?5����W�}�W�}�W�}�׶���O����x��ǯx|"��H�S��ί���N�M����M���k?��y��<~�����<��~�s���ke�����O~��W�~u�W�~u�qE��չ_�ȯ���<>�W��L�~m�:�+j����`��C������k?����
�@�
�@��O~m�j�������|C�G���_���S�*د��*دe�W�~E�W�~-#���_����_m�D����~�M���+D�B�+1��'���_�Հ_�����O~��W�}u�W�}�,���۾��۾"�+Ҿ"�+Ҿ��+����[�ͯH����"�ʯ���j����j����W~}���b󫵾Z뫵�Z�+����k������u>���g&���Z_���G_}��G_}�Dޯ?�O0��x�֌_��9_��=~�S>O�!���|���|�2�+s�2�ke��9O��vɜ���Zl~���Cb�+��b�k���4_��'�2�+s����D�<���qE}��W}��W}��W}�,���_�ǯ��ZF>���1�����+��*�+���諏���xy}�m���d��)>��N񫢾��+����裏5�WE}U�WE}U��N�k���Z_;ů��Z ~��WX}��WX}-�*ꫢ���k��UQ_�¯���~U�WE}����|��!��f|"�s���j�������dz"���G_1�m����W}�'���+����+���諏���8�>�꣯>z"��x�LO�!����<��U�W2}m1�b�{�rb�|�2�+s�2�|C>1�����b~%�W2=��w�I����WE}�:�*ꫢ�֟_a�V_�����꣯����|6�_ѯ��W~}��Wk}��WX}��ג�k��V_�ͯd�B�gz�ί}F�h��Wl��a�"��,�"�;�^t�~?��+�>޽�+�>˽�C�N��н��H{Qy���f�"�;�^����r/�S�E�w~��C�>�=~�!~Gڋ|ۿn/�=����)_�{�}�{������"����"O�;_�Qg�<��{��������y����y����"o��x|���}T|���}T|���}z|���c��>*����_Ĺ��/���_����yE�*�/��U
�_���C�Z�y�ߏ�/�\Q�����C�Z��	��"��x���E���'�y�߇�y8�����C��"��Ĺ��{����ys����"��,��� �yEg!��/��4���|yG��E\��"j�A�/�����ƽG���s�~�}�W���
/�N8�hj�w�)�`�Wt���_�!|�����s9��/��|T��ȷ�ù���r~������w2��'r�P���?���Ї-:��Z�o��D�/��$�E^��Ao���"%�/������;6�E���7�E���p�q'hD�W��6]�/���>��b>���§������KC��_����'���<�O
�y.�!��_���N���<���^�Q}�@���C��~���ț�)j�_乜Ԍ�ȷ�������G�O�c=�/���_��ӄ�����C[�����u�"��P��O��s(�~����1�/���(��w�~[��~��r�l��E�����"�蜠@�E�	�	n�E�{G"�E^��A���9~�y�E���yk�"NO���|y��/�~a�'���E�� E�"~(�y?@�_�!0��ה�}�G��+:shE���Š��E���E�"�N��<�s�:��Z�	|�|��	��<�����y.�	����x.�	u�/⵨�~�U������~�
�y���/�\�!��_ď��
h<��+P���!���|y��E���� V���;s��/�~���~���9��_��y���E^���~�w��V��y.�"�E���~�Gu�ё�"_�1T��_乜L ��7��"_��~wE�"_ޡ��~�G���8P�/���=&��E�Gj��/�Μ�C��E�i��~e\^�i��~�Wt�`�_�0�����9����~�Gu��'r怴_�QC�1tC�1��~ui���>t|���s�9���W����~�/���CФ�"��>l!�_�����WtR��"�c;a�/���r����Z���NL��<����yT�(�E��H�����C>��z|�ȗw���"�:�(�~���a��rP�y�L����_�f���������Em�D>�a�_�!|p����+rs��/����A�/�L��W���Ad���;�h�~�W��8�p�/�=:�p�/�>�!�_��u7��/��"���z�%�/���Bd��s9�@�/�>�Q��"�専r�ȗ�����?���v~��_�!V �y��/��/:�_��	������	�?��Gm��~����?
�_�����ݟ����E�<��rb���F��O����?��_�Q��,�Ӏ��O��Q��"����ysxp�ߟ���rO�O���ѷ�"�,�ߟ���m��O���c�}"�O����?��'��ٟ���_��|y��'���՟��V�ꏆ�y.F����V��OX�	�?a�D�����SQ*�OE����"~ڟSNk�i�?��D�8>����_��Ok�i�?��_�k9�h�o��E5��|�<�}��O~�i�?��D�	~U�ɯ?��D��G����_<�}����C�{�O��ɯ?��'���C�\��O�"��s�'���'�/��ZZ�Ok�Q �"�E�������V�ꏶ���r�)'����3�|�+z�_���H�V��OX�I�?z�_�}�Z>-G��/��L��j�y0�ȗw���'���%���C8`�F��Q3�"��̡��E�/~q�)�?
�_�k9Mt�m�/�9�t۟n��mOč���ɤ����e��kE|-���Sw��/�&��O�=7G���?:�_��0��O������9G�=���C?����OC4���s9��1D��<�3G<���?�'��t�y.~]�ɯ?��_����SQ*�j����"�6=�/�=��"A����#��/�N ��'��h����D��I�?)�'����5�/�\�����yT��/�\�
�_�0J�|�N��'���,�����O>�?Z7$����r��"�O0�ț�Hӓ��<��>�y�菗�N8����/�=:�����Q��"�=��/�
�?�'r��P����?z�_��N�}"���B��yz'���S����yW�_B�O��	�?!�G�����#���y�|�����Ou�Q��"ߐÊ��yTg�6�Ӧ���yɴ�6�Ӧ�̡��E��3G��	�?!�'D���=�/���hm��M���6��B�Ou���?j�_��E������+�ѭVr������L��z��k�e�n�H22�IDeD�����B�+Ɇ-a��qԔ�5gk}�ߨ��zEf��E�}�`���A�| �����MH��$��9҆��J<m����䃤� )>H��⃤� )�O��Т!-��xD�>�6�X� �������pD���f�l� �>��J�j7��@4�+a&�B�P�@4�+q�!���4� ?H����� ��Ag"�>ȹr{K<"$r�@��+q&�r���_�O"�>Ȧ��l� �>�"�-���LD�y�Ax| @��xq�F�|�'o����<� <���㯄#�'o	����W��1D���_���1�T�'%���E�|1�%~<���� b>��"惈�@>���i�f���W⸸$u>m��yK�,VVD�ǡ3!f��xB��C�"u>H����/�毐{V#%�.G6}�'��y�A�| y��x��4��<�@��+�҈�Č�&� � b>��J<"�4���&� � b>��J�xVV����A�| @��xD:�_�SHB4�+q&hC�%�6m� � �>��� � u>������@�+q��L�o�6D�|1�o��A�{ ��%�R�_�O� �=�r��An;����A�;�m���sr�-��Q�!� k���u���A>:�G�� �b)� ��� s0�:�4㩃 s0x:�4�� ��[���=�`�ts2�A�9)��FJ��`�t���A:�9#���s�|FJa� $�[��3?:�̏��A�9�4�� �d��Ls`��d��Y�� s0,:���r0?:��a�A�9H+â� sM��A9��`�s��9A� (��[�|�sH�����-q������4f>�� t��[�L�C��4� t$��8q0�9H��A`)��B�����`�s�V����� �����r�V�@c�� s`��hCA7aNs:�49���,}	�8�Xw�� t����q'��A�8�c���q�0�A�8H����q�0��-�b0�`����qK	�`�t_/<"��r�CB��H� ��?�>�H� �IS t���đ,W��@�8H	� a$���q0��%�&hC䐃r�Cr�A�%~<&i0����q0�9��� ;�in�G�L�8�W-	� ;�~9ū��pR�A8��D��pK<"/d�-q�����A�7�ġr�x�2�9����(^��v��n0͹%��� �$y��n���A 7��� jDm���Q\w�m�O� j�j���AԶ%�#}��m���A�6��o[��@n�&C�� ��2�A �%�nB�6�L�f>�ۖxDV
Dm��m���AԶ%��D 7���^vpt&ҷA�6��#���m0,:�n�3�M�IgbXt���E�� ��o��m0,:H�3�������xD:����n�b��H� �$y[�L��GI� �r��m�r�A�6���?�u�ۖ0��k2�AF7���� D�O�nB�6��xn��J�!�r�@n��A 7���`XtK*m������`�s��2�AF7=��m��m�O�`�s0�9�¶�?$�N�,l|m	C�,1��Y� ���A<�%��>A<6�Ƕġ�'H��� L��Ab6�Ƕďg���� da�,l����A6�x<Ӝ�xl���A6��_[��� �HR�A�5���\�A�A�5�DZ[� H�)�`jr�rR�A~5��DZ�HkK=��djCF$󐃰j�92�A�4��� :�D��h0�8���k���-�X)�&Ҥ���``q�9r�A(4�Ӊ��g0�8E�"F����h��At4EDG���A4H�AΖ0T�������Y���vC��lgK=�	�A�32�=[�Y� �s��Ph
���� ��A�%N�Ph
�A4H���[�hCL'F��`q0w8H��$G�LЬ����`:q�&�[�P�r�����``qi"���``q0�8��� ��\��k>����k2�8	����A$Y�$�da���I<6k�ǅ��$D��h�I�I�6��&Ï���I�6��&�[��I�6��&!�$D�LN&
'Q�d�p2Q�%~p�$��,-2��o��m�M�'�ۖxD8S�M�������I 7	�&Q�$j��j�\m2d82�Dm��m��Mr��D�$W����$W�LN��IԶ%�C 7�;�dt��n��m�O7!}��
N��ɬ�$}��o��m2>8���o�\m��MF�&#�\m��Mr��|�$W��!�Q�|�$���E�b�o��M2��0�$���v�a�Il7	�&��$��rs�@J��`��8��ܖ0� '��d�o�M�I 7	�&��$}��o��m�M��I�6��&Q�$D�$f�)�-�,j��&������`�d0pK*6���nK*-���I�7��&s�[�X�Q��(�$����Q�I*8I'y�$�LN"�-���rA�#���3Xn��M�#(���Tp�
N�'A�$(���Tp�
N�'s��Tp�
NR�I*8X���[�i3�8�'���H�#	�$a�ĉ3i|�0N��I�8�a�$���q�0N�'��$a�$���q�0N�I�8I'	�d�p�
NR�-q�\�n��b�E¸%��6����19I+�O���u$��hrMN�'i�d�q2�8�t��5΢)MN'i�$������r�VN��IZ9�!'C��hr2>�%��J�r'��D��hrMN&
'i�$��n���j�Ls�iN��IZ9�;���u1�$朌"Nb�I�9�;�$����I:�(�$���sK<"x�"N�����$�䣓|t��N��ę����Jd:�L'��$2�D����I>:�G'��$�L'N��ݗGd�C�:�L'��d`q��N"���d�q2�8	V'��$X���`uK��i�D���I�:IQ')�$��H/$2�䣓|t��N&'���I�9�r��`u2�8�L'��d`q�N')�$E������I�:�L'��$2�䣓��I>:�t�䣓|t2�8�t�L:N��I��%�����jn��-���IH;	i'!�$������v�N���<�drK�x���xD�Q�x��'��w��Nf+'��$ݝ���tw��Nr�In;���䶓�v2[9�r��G��N&0'��d�r2[9������w�N�-��Ӧ�2���*}�<y��<�y�$O�RN�&'��$)�$œx�O2�Ɉ�$���(wK�x!��c�q2�8�r'c��(w��Nr�In;�m'��xڬ�Hw'Q�d�q��n���u�nI����09����E�!<��6���$b�RNR�I�<	�'#���Ɉ�$O�$œy�IR<I�'�[�#���'Ï������$b��CN"����xD�С1�8I�'��$u��0Nf�a5D6=ɦ'c��lz2ø%��F\=	�'��$u��Γ���X�d�q�MO���t�8�4���t�$��dӓ�y2�8��'�<,D�N�L'N�����dq2w�%��zK8"	��0L'Nr�I�=�N�$ؓ{�`��j��sH�'	�$��$ؓ zK�,�C���yO��yy�O��Ix<	�'��$)���Y�ɬ�$𝤻[�	�� ���tw��N��-q\,1Hw'��$ݝ��[�qq�h
䶓Q�En����c�.��E���rQ�"�]��[⸰�*r�EH�i�$��|�M��v�.F$��A�`��v15��m�ĹǢ��\�[.2�E��%~<��%�#*�")^$ŋXx/�-q�"���V$�[�aiER�H�I�")^$ŋ�x�/b�E,���\$ŋ	�ER��\d��x�.)������tw��.��E���rQ�"�]����-�g�'G���r��s���.�E���\R.��E����\�V.2�5�9�q�Ÿ�"<^$�[⸰;\d��x�/�E�%��tw��n��=�bs1���r��b�r�.��Ÿ�"�]L`.�E����\���q�E���rS���v��.F$��"~]L:.&!�b�q��.B�Ť�"k]d���u��.��Eֺ�Z�ę����.R��l�b�r�.����"k]d��uK݄q�E��V��"]A� ]���y����u��.��E>��G#���s�|n	�J��k\���hrM.r�E��[� x!'.��-�y!:.B�E踘t\���p.���s�ݝ��-q\���A�x�,�� �������EP�
�"\D��p��-����EP�%���p1鸈�ġr�@¸%�����6A����#n���*�I�E¸~\?.B�E踘���Z�H	�"a\ĉ�8q'.��=R�>A¸���br�m�HS �[�{�po1��Ï��o�-b�El���Ï��n�-�I�"�[$y��n1鸘t\�v��nK<"�I�Ť�"�[�}�zḸ|�\>��-��E��H���"�[dt��n1�������n�-2����"}[�o��m1�����"�[r�@n�m��P��IF�%��f���b�q�-½-�t&b�El��t\�v�I�El�����@n��-�E<��;\_��ki-"�E~�ȯ��"�Z�W��jK��<G�i�"MZDG��h1�\L�4i�&-��EN�%�2iҖxD��	�i�"MZ�D��h�-r�EN��	�"�?��(9іp��zb�xؼ�E\�".��t�"sZdN���E�������Ŭ�bVpm: �����E�����[�y�߼��&-ҤE���	�"�?�@�%9"���b��"�Yd;�lg1+��{��"���H`
p��,��Ŭ�"�Y�
n	�`|p
-B�E(�H�q�b|p1>�H�	�"Z�=�!�Eܳ2\$@[��s�ph$@�h� -�	�"Z$@[� h0,.���"Z$@���-��}LB�E(�E\�D��hK<mV0�D��h�-r�Ť�":ZL:.Ҥ���"`ZL������b�q�L-�a�"�Z$S[�h��U��jV-f+�պ�G"�E������"���Z"�E���\e."�E~�ȯ�ՖxD��墌�j]:&��	�E����	�E���㖋q�Eb��\����"[�c�xl1[�H̶�ɡ�2n���GO_%�[r�����"�[R.��E���!�"�Z?.���ϢY�-B����"W;	�NB��Ɠ��$�:��N"��H�$�:��NFOR����$�:��NFOR����$�:	���#�s&3�[� `C��kK�1M���,�$;��N���ɓ,�$;�<�<I�N����-q\��I�v����Vn�GD�7	�NB���$D;	Ѷę��M�-Or��\�$W�ǅ�n����i�e�L`�r'�ۖxDz!��P�IFw�m	G��&s�'I�Ilw۝�v'�'�ݖxD�*C�[� �D�'�I�w{'����I�w��dt[��i|�j'C�'Q��P��P��P�I wȝr'��I wȝ���P�8�����8�/½�$�d(�$��Ag"�;	�N½�p�$�;	�N½�p�$��������
��|���[��rL��ĉ'��'	�I�x�0�L��$�'��'��'9�8���I�x2,z�C���D�'â'��I�x�0n�O{d��$�<��<��<�&O�ɓh�$a<��?��I�x�0�$�g�.d��d��$���E_e��$�<�<�4O<O2͓iΓh�$�<�&Or�-a\D�'C�'C�[�L0�y2�y�i��[��g�`�4O2͓��-���h0L`�$�'��[�iĜ'1�I�ys�R�Ĝ'1��Y��H>ϤO$��[�h�i���'����I�z���L`��V��[�YF%�|į'��I�z&��Z��&��'!�IH{�n	Gdt�$�=�rO�ܓ(�$�=�mOr�-q�t&rۓ��$�=�=�'��E��%�W�E�c~�$>��O�-��~$�=	|Oߓ)ӓ�$>�E=��OfQO��X�$>=	|Oߓ��d��d~�$>=��O�GO�GO�EO&CO��-q�阤�'y�ɰ�I�|�'���L��L��$�'3�'I�IR|����'�I|2�y2�y��x���'I�IR|���'c�'I��d�894�I�#<>	��ď��1z1�D�'�I|N��������xBt&"擙ϓ��$b>ɓ��A�J#O>	���xD:��Ix|�$�'I����x�4+�@O�@O"擈�d�$<>I�O�9O�4���bt�dN�$b>��O�2��)$���Ebt�dt�$�>�<	���?��,H��[�	�)%A��l��l�xB���<ɹ��#�s��Or�$�>�ɓ��dD�$�ޖÏ��j��HnI>���҇�ɓ�ɓ4�$?I�O���-ɸ�+d�Df�%�e1�I��%���Lb���dN�dN�$F?��Ob���$F?��O2���d(�$F?�<I�O���d�dt�$Y?��O�	̓��d(sK*m��d(�d(sK͊H�$�?��O���q˓��d�$�?��O"���̓�̓��$�?I�O"�s����Of+O"��H�$�?��<��O"����$l?���CS F��J��%���$ ?	ȷď����H���'���<�I~���D�'��I�}j�L:���[�9�/wr�P�$�>��O&��)��N�}�s���[⸸D"�>��O����$�>��O����$�>ɹOr{��xD	�I6�%�6��I}�:���{}��b����0z"擩ɓ��$u>I�OR�AʓAʓAʓ �$u>����#ҙȓO��-�㹇Lx|2�y�$�'�I�{���'��I�{ҞR�LM�LM���'��� �I�{2H�%���@,|2[y2Hy2Hy�'���[�X���$���� �E|�oI����_��H�/����"ݽ�a�?��"��N��N�|/ߋ��"ݽHw/��-�(D���En{�^į��Xį[��:Yį3�����EH{�^$���E�z�^���E�z��^����)�8����"2��G���(1c�)�E�z�^D�Ï)��X�Edz��^���xD<ZD���Edz15y��^LM^�[��Q�,)�ġ������"���������m/rۋ�ʋ(�b��b��b��"�|/ߋqˋ�wK�(�"ʽ�r/�܋(�"����g��E�z�^��)�E�z��^��WЬH>/�ϋ�rK��E4y1�x1�x^�A�E*�%�&�a�
/�/�Ë��";��/�T�"�� /�/R���Ë��"(�
//�Ë��";�
/R��pK<"V:��"�� /"�-�M�a�
�ď����Hb�c'^ĉq�Ev�%�yȋ��"N�����fj�"a���r���"a�H/Ƌ8qK<!V
������E¸%~C\�0^I�a�rK<!z��8pȋ��"a�H/Ƌ8qK�x���/�2/��+��[�|�:H/R��TpK˂���^d�A�EPx^��Ex^�}y�E�w��]�}��W�M���.½�ϋ$�bt�"���ȥyߖ8z�E�w��]$yI��4����a�bt�btsKrD�6=���"���.�-񄸕BFw��]dt�U܃a�"�����.f>/f>/2���ϋ�ϋ$�"ɻ�H�.���$�b��"ܻ�.b����"������.��-�hC�o�ӜפM�9dt�E�v��m���M�>�|n��Mgb��"����M½�p�"ܻ�.½�poK��p�"ɻH�.�@��s���]$yI�Elw�]�vc�I�Elw�]L�^$y�����d�E�w��]L�^D��Ex^�}I�E�w��]$yI��,��m3��%��E�w1��%�*͊��b<�b<�"�� /"���"�� ��#ҙ�~�H/½-��i0̵^�{���\��\�8:A�E�w��]$yI�E�w��]̵^$y�EFw��]��^dt�E �gG$}�>ksQF�v��]�o��E�v�]��A��%��!2�����4��@�b�uK���b�uK<"݄��"���.򾋼�"�H�.�����bl�"����.�f/���$�"���.�f/ҷ���"}�H߶�Ӧ�lzΦ��m��b5D�wm�զY��]��^D����E�w1\�%��ڋ�pK8m�Ë��b�"N������q�f"a�H/Ƌ��-q\2�{�C^�S���Ey1��%�.G�x�n���
�b��"t����/�ċ8�"(�
/���"(�
/½�!֋p�"ܻO��.½��Ջ��"���.�)Ӌ$�"����� ɻ��.<����%JFw��]��
â��El�%��;��^�n���Ͱ�E�w1,z��]�}�[⸸j"(��2�)�)��/�ċ8�"N����qљ)��?�C�x�0^ĉq�Evx�^�}[�g�:� /�@�ֱ� ��׏o����_ ���&(�IoR��T�f~�~PblFJoFJo�-q\�M�x3ez:�L��L���79�My�Cބ�7���H����������My:����7â7���d�My3z3z�C��79�My:ބ�7c�7c�7c�7i�����D�7��������M4yM�D�[�	��ك�Dy�Cތn�D�7��M4y3�y�C��i��in�OK#����I+o�ʛ��&��I+o�ʛ��&a�Io�-��srhVLs�d�7A�MPx�
ޤ�7��M*x3z��7��M*x3z3zn�?&l+����s=�iΛ��ft�&N���IoƛiΛ��&a�Io��-����Io�-oB�-a������&orț�fDrK�xz#�7#�7#�7#�7�����Mz�ބ�7S�[�PiCRޤ�7)�Xn�՛�&E�IQo)o"�-�4+"�-�iC�7a�Mz��LM�$�7��89t&�Л0�&��u�&���&���5)�M�z3ny3ny���d�[��~$~��_o��-a\į7�����xDz!��[�i���d�w��_o�כ�ϛD�&~���E�z���x�įwҬ�_o�כϛϛ��&��	i�ˑ�ބ�7Y�M�z����7��[�ǳ�"k��HKc��&~���ݼIdoٛD�ft�&��	ioBڛ��&���Ido�9oBڛ��-�'G�z3n�%|�$�7��0�$�7����M�z35y35y��n������į7��M�z��į7�7���l�M"{���$�7��7!��l�Mn{���L`��7C�7!��P��P�xD�����M�{���[� X1[�%~<-�(�&�������ro&0�į�eQ�M�{��D�7Q�M��%���M�{��ތnތn�d�7�M|��Ls�Ls�eޤ�[�	�	|o�ܛq˛q˛(�&���H�#���E�#ݽIwo�ݛt�f��f��&�	|oߛ��-ɿ��Yl1�y3��%~��m�כ��&~��_o)o�כ�uK=˨I"~�N{�`���fD�fD�&E�IQ���|tK�,^��C��C�D�7��͈�M�z��ޤ�[�i�@"X�	Vo�-o�֛��&k��Z����`�Zo�֛�uK�x�Y�M�z3[y���d�7Y�M�z����V�d�7��[�ǳ�!X�IQo�!o�!o�֛��&k�����_o�כyț��f�frK��09�H��7��Mn{��ބ�7!�xD.�6��t�&ݽIwo�ݛt�&ݽ������	|o�ܛ�vK�,���M�{��ޤ�[�i�b�&�����O��4��-��/rۛ��f�f�&ݽ���Iwo�-oߛ�w+���&�ɀo2���&�ɀoߛt�f��&�	|oߛ��&��>�(wK8!�ݛt�&ݽ�_o�כ`�&E��E�a��&k�IQ��#��b��&k�����_of>��q�s����â7��Ͱ�M�{���7��M��%�%S�[⸸�,�Mx|��L��d�7c�73�73�7�����8.�_�7��8z�[���p���7c�[� ���2���&)���	�o��X�&�ɀo2��xK<!z��M�{���į7s�7��M�z��į7��M�z���7�7Y����M��%�*/dRԛ�f�f��&k��Zo�-o��-qr�;��C"���>$�[����C"���NtW+<"��C"���>$���C���n��S8$���C��0�%�p�Z�և��-�XRԇ�-�q�?�V>��#�[⸰�8�i�8_�ܻ��g��?������C�%N!��!t|HƇIǇ��a��!t|�t|�!rȇ��!N|��Ç�ŇQć��!(|
F��Ç�Ç8�!N|�F��ć8�!N|����-q���Ç��8����ć��qK�UZ��C��:>����C�%����!t|J��8�c���pD��-a&H+��'hCAbrK�j�!�-��iC�[� X)M>e>��i�CZ��V>D�9�C��:>$�	����C��%~<����!a|H��s��Cn�MKc��a��!�|��|0̇ �a��!�|�|�9��q��.G���i>d������C���i>d�i�C4�M>����4�C���0>$�	�C���0>x>x>x>D���C4�M>D�9�C�%��^�t���1,�`>��C��%�+>FJ2͇ �!�|0̇ �!���;��)Ӈ)Ӈ)Ӈ��Iz!��Ô�C�%�^�,�C��n����%-���!���J�"�|�9��A��9b·YԇL�a��a��!�|H>O�χL�!�|)}0�ġ�J+�#�#�O�s�42͇L�!�|�42͇�чLsK�C[�9�C��C>�#����H��H�S�rȇ��!t|Ƈ��!a|}}H��b5D��:>̏>�9�C�0R��C>$�	�p�$�	�C���0>�A�C*��
>��Ϥ�>��>��>��>$�	��H�ð�C��'>̏>̏>$�	�C��0,�'>d���C*�0�>x>x>�<f>�ć8�a��!;|��@�@�$G��Hg"N|��ćχ�͇8�!;|��|���o�i·��!a|��|��|�!f>���a�!�|}0̇1Ї1ЇL�!�|��|H+�ʇ��!�|�&rȇ�!a|H�Ç��a�sKrD��X-VC�[��9�����[eQC�'>�nn�Ϣ�i·��Y,jf>rȇ�-��L��i�C4�:>����C��0���0n	O���0>ĉq�C��0�%����:>ĉq�C���>d�A�CP�0,��>�>�n��b�D���0>d����d�C��'>�>�fŰ�8���}�EBǇ��a~�!�|�!�-�iiĉq�Cv��>d���C*�0��>�}y�C����=xn	��4�C*�%��!|� <�9��A�@b�sK�j	�ġr5w�rL�>�|>��i�C4�M>��n��E�"�|�&�ɇh�a2�!�|�!rȇ��!t�ϑ�D��0R�:>����Cv��>L�>d�S�#�q��H��H�C��:>$�	��,����8�_D�����,�C��0n	�E��:>����8�9�è�xD�ץ`>��8.Vi��>$������8T���x�4+�Z��b����C>���>L�>L�>L�>L�>̵>d�)�xDZ��C��0���>�[�h|į[� X�]�#��Q�Cn�0��>D�[���L���mrۇ��!�}��}�m_r�-��/Q��p�K����D�/Q�K��%~<��d�/Y��Y��������K"�%�%�eF�%�}�__�Z����\�Z_&V_rۗ!֗(w�1yDLK�/TV�X�e��e��%<~u}	�_�㗤�e��%<~	�w��A�s.�K��2�2�D�ľd�[� ݄Y�w����/���H�K����̏�d�/�[��� ��/�K�2?�%�6/wb�-q\(j.��K,�2x�%���%~��_�L_�L_�L_��<�%O~�2��H�`��%)~��_b�X�%~��_2��xK6�/��K,��d�[⸰(���n��BӋ�#�����pB�/��[��ɀ_2���ӗ(�%�}	i_Bڗ��e~�%~�k2�!}���e��e�sK*�mRԗ�%2}�L_"ӗ|�%}	C_�З��%�|I>_�ϗiΗ����I>_b�-�ym3���|�$�/Ӝ/Ӝ/���4�K>�2�����n��i��i��/��K�������/)�K��s�Ĝ/�/��K���|�$�[�h0��[��&L`���/�/�K��`��/9�K��C�I�!t|	_Ɨ��e��%N|�_��-��&I7!t|���H�!�|�!_BǗ��e��%t|	_BǗq˗q˗hrK�I_�-_BǗq˗q˗h�-^[�Py�3[�:�R�ĉ/q�K��'�L:��5��5�$�/q�Kv���/A�K*�2��2�����/y�K��2Q�2Q���$y/I�K�����
�dt/��/������`�K����$y/�}/��Kl�2����m	�8yw���Ƚr/����ߖ8z^�r/��K �Ƚr/�}/�}/�K �ȽL�r/cz[�9r���%�{��Ĺ�L:�亃poK=�� _"��pK�"�6Đ�xD��/����K��ѽ�j/��K��.�S�/!�K�����h[¬.��L��o[�Pi0r/C�/C�/�K�����������r/��������Kl�۽�v/�K �Ƚn��31+�%�6D����L�����@l�%~����eV�%�{��^2����%�{	�^�__2�)�\Q۽��v���R�L����v/��Kl�۽�
�L��v/��Kl�2��佌��$y/I�K��۽�v/��/I�K���佌��{/��/y�K��{/���m����$��O��E�b��%�{I�^b��������$�M��H�#�{��Y����t9½�p�%���	R��Ь͊a�o�%~=���%}{��^r����%1{��{	�^B�o�%���6��K���_��W/st/��K��2G��r�DZ/��K��24�2!�2���_���$S_���^b���%�z��^��^2����%sz���d�0_̾�$S_�A2��L�$S/��K�}�O�Gd=A�C��I/��KN�}��e���%�est/���h�w�����%szɜ^2����%s��PQ� ��a��e��%�zI�^��r��b����e��%szɜ^����%`z�|ɜ�75J��K�#s�Z$z!�/����O�_푉������)���Ѫ_-E+іh[�Cm�1������Î!�r�����7��B��r��;�W�9H����M9ߔ��|^�y����2WS�cʘ�w�yL˒�[2�%cY2[�m�1�c˹m9�-�q�G�{�G���q���c\��+su�Z�2W�rm,��!>4�����x�!���S�hC�18�C�j�_�!>��l����x�/Y���1�s�x�����_MƗ2>�^��d|%s_2f�v��d��?����X��x���uC������|���c���s����u?���ɹ���z��d���~q�������!�6�׆�Z�_��M!�KY�j��
��B�)�n
����~59��Z���xXH-�k?x���Z��
��B�*�_B������Rs�xS����&ǐZ*��
��B|(�́�W!����̕xI���xIH-�!���x��̳�F���4)��H�:'��I��H�_�G��Aʵ�RӤ\�)�y�5�R���/)�Kʵ�r��/)�JJ��R��xD�5�rM��)�yJ�r�璿��7��H��Sꈔ5SJ�r�\�)�y�u��fJ�-R��!�fH�?H�uO�G���RRo��A���%k���P�G��%�E����%^R�%%�EI}P�%�Qr�\�%�~ɵ_R3��AI}PR��SJ|�d�R�%�@�}�d�Q�%%~P�%~P�%~P�%�~ɵ_��(�J�UJj��(�k)񈒵F�Z��K���ߘ�S|cJ�1�ޘ�/S�e��L�)5Ȕ�b�GLYCL�#���?��^�R3L���Ɣ5Ĕ��)~0e1�#�x���Ro��z��|R�L�A��˔d�b��L�)5Ȕu�/����RGL�)^�w����xɔd��L�)5�/��%S�d��,Y�,�%����K�`�:e�G,�A�� K�-�K��˒dI�ć��K|c�o,�7��ƒzcI���K�xɒ��%^��K����kI��d�aI�dt�o,Y�,�%���VY�K�%u�/Y�K|cI]�dM����K�`�lY�l�-�Ɩ�b��Ɩzc�ol�#�xɖ}�-^��K�x�/��lg��l�-���_��*[�A��/[<g�>Ȗ�f�m�K�����R�l�-k�-5Ȗd��l�-���_��%?�����I��ee�m�-�-�g��Ֆ�Ֆzh��m�-~�ů��Ֆ�gK����zh��m�#~uį��9G�#�v��9�>:�aGj�#~uį�xΑ}�#�s�s��/G<爿�#u�9��r��9R��s��Ց�爇�#v�Î���<�=�WG�LG�#v�Î�HG|툯�#�v�׎x�:�CG|�Y����x�o:�CG|�Y��!�Î�aWj�+~uś�xӕ��_]�+�t����WWj�+���R7]�+�CW���Z��~�����t�6�R�]��+>ye��O^Y^��+>y�'���O��W<��z��'^��������Wj�+>y��x����W֗W<�J�w����W�+>y�'�����+�x�^���}�;�����R�]��+{Z׼�k�V1�!��x�C����'��u��y�<�u�5a�[�w>�knM�B�k�!��x�C��!L�&z<��!��x艭���'�0ѭ������q;=��nM���qOݚ���9���]ᮇp���ᮇp�C����c�C��g᳇����ڹ5�t�=֧C��!l��{�=��nM�_��x���a�[��Ћ�0�Cx�!���{ֶCx��8�!�=Xa�[�w.��V|+>��!>.\x�̋����5��|S>�)C|\8�1�ǅ=�̇p�C��!��~|?>��!��!� aʇ0�C��1��)��O�+�,Lyk2���C�Y�������̇p�C��1�c�x���|��C8�1�w�)aʇ0�m<F�O�x����!��M��yV|+��E�!�|ޚ�E�E���va����C��r��=���qḇ0�#�:�����q���<�:��B�}�p�C���d|\���>�V|�����#��
��0�C����m�s �yk����Ix�!��μ59��H)5R���P��W�!<�}��C£���W�!<zkr\�aχ��C��!��H��u&�}��9�Q¨a�G��%�M�&��憰�CX�!,�H�5��[�yK�+�ۇ��CX�!,�H�iR|-��R<L�����^~/?����aㇰ�C���8W������C����o�ׄ��e���xXI�$l�6~�K!9�xX��	?J<�Ȓ�_+Y�	C?����a�GImV�k����G�����J�NX�Q�V�~?����C|��ׄ���a�G��	�?����a�0�C��!L~/�e,R���UIm&��vL�0��p�C8��x\a�0�CX�1�9����MS�+��ǔ����5ν0�C��1�7�����CX�!���R7	?�������o&�?�x�p�C8�!����M��)����C��!�~k2/RsM�0���0�C�!<���ߚ���M���&�+�C��%�#��v,�����ߚ�E<Gx�!<�v�?��A-�&�����Cx�����,�%5ג�k��I�@k2f����`,���g`,�D��30�����hM�+~%=�ɼ��,Y�I/��^���s�?`H/��^����C�0�`,�%���YRIo��ނ�d,�W�[0��`Ho���W[|h�I��>�!}c��Io��ނ!�C����a[�+�[<l�_m�+��3КC|H����Ln�7I���ނ!}C�ƖI�ƖIz����0�?`H����!� C��!��ز��?����a�[��ٲ���/��a������Gja��ƿ5��/��?��������q��:�C�G0���5��MG�!�-�[0�xΑ��#��#{��G0�?`H����!�C�Ƒ�GzZ������`Ho��ނ!}C����G����M�0�?`H/�8�aG�&��0��ߎ�C��a�Ǒ�H=$���\�+a��o��M��a��0��7]�!��[��!����?��W������Cx�!���R��?��Wja��oN�?���p�C��q�_������Ǖ�!��p�C��!\��R#	k?���Џ+�+^"�^~\�~��­�dt���!�!|{<���p!|{�����¼�0�!�{���¼�0�!�{�²���!�߭���9���X�d��0�!}k2fp�!,{�£���!<zH6x{�0�!�xk�}�V	a�CX�.<���C����.<��a�C��\[���!|v����]�p�!�uHFwkr\��C��>;��a�CX���>;���C��>;���C��;$�5�x�p�!�v��]��,���C��|��:��nM����;$�;��nM慵THx��l�0ۭ�X����a�C���:��nM�W�Or�[����-�َ��D�C��C�퐼����l����{��C2�C��<$/<�����CX�.�5��a�䊇d��&���`H�xH�x�£���!�ykr��Bj3��oM�Y|M�F=�Ga�C���<�3��C8��<�)����,�&&Lyk2��k�0�!xH&y�I���M����)a�C��9�x���!�x?ޚW�I8��<��<$㼭N��}���5��[�㊿S���!�xH�ykr\���3a�C���<�)a�C���<�)a�C���<�)a�CX�V<�oM�!�TJ-%\x��{���!�wk��ޭ�牿����ݭ�yH�$lwH�y�ݥ�d����!�w��q�p�!w�%k:�=a�C8�f;���C��>�59_��Qa�C8�l�����q�p�!w����v�&�/��>;��a�Cr�CX��5����!9�!�vH�z��q�䨷&c���&y�����xݔ�������d,�k�����&�_������^2�q���a�C�<�a�Cx���59��H�q�Q�M�!�C����<į�x�o�;$��59��>�v�䷇��!��!�wH�{�0�q,�0��;�;$�=�o��+xޚW<GX�.�5�x���!�x�p�����$>��a�C��Cx��;$�5�x��ݭ��+~��6�,��<�.�5��a�dɇ0�!�xk2WR�-�%�'9�!�y{���ɘ�'�x����X��=a�C2�CX���~<�a�CX�V<�a�Cr�C��~<�a�C2�C��~�5�+�5ɦa�C���<�)a�[��C<Q��\���|e�\8��<$�>�3�-�&LyH^}k2�:a�c��	S�/�ߚ|��&�/����<�3��[�q��R�dɇdɇ��!<zg�%�dɇ0��1�s���C����|�s�ɡ�#�#Lyk2�!a�C������<�=ɵ��C2�C8��<�3��Cr�C�<$K>$K>���C��[�s��J2�C����5��R�9�9£���!�yk2>�Dɫɫɫa�CX��=�e��[���W·���!y�!|{k���C��n=�[a�C���ܤ��=�ea�C2�C�����kW|MX����=$�>�ya�C���l��59��f·�dη&�"�$�>��a�C��6>��a�C��6�5�{�D��Cx�����d�'%�>$s>$_>��ɍχ����ߧ��)�}
W��էp�)��)��)�}k�]��˧��)�}
��ߧp�)\}
W��%����ڧp�)}
C��Ч0�)�|J�|
C��C��է�Ч�Ч��)9�)��)�~
���9��9��9������)<
ϟ�%ߚ��z)��)Y�)� )� )Y�)y�)�
�ߚ�/���?��OɃOɃo��+�k�p�)��!~%�~
����0�)�}
k��ڧ��)�}
kߚ�k�����>��Oa�S��Sr�S���>%�<��O��S���d�K��oM�ǚ+��O��S2�S�����>%�<��O��Sx�^>%�<%ϼ59�x���)\}
Cߚ|�\K���)��)�|
�¼�0��1�sB<G��6>%=�yO�BO��S���=�yO�GOa�S���=%=�k���59���d��p�)�zk�I�%���¨�d��&��F=�GO��Sr�Sx��#$�59�xDȵ/Ly
S��d���sK���S��V<%�5�Gʵ/Ly
S��䔧䔧��)��ɘ�7�QOa�S8�<�<�=�=Oa�S���<�)Oa�[���uO�o��*¨�0�)�z
��)��R������)�y
g��p��X�V�<�=O�$oM>Oj��S2�S2�S��L�L�=�GO�$Oa�[�1�=O��K��!<zJ�xJ�x
���5��5����)�yJ�xJ�x
�ޚ��xNI]"�y
g��ޚ|�/%�R�/¨�䏧d��0�)<zkr\�i�QOa�Sx�,�a�S��S��<�3oM�����<�=O�O�Oa���#��n=%W<�Qo�Ǖ\�=�=Oa�S8�~<�O��S��S�<�oM�,�3e-$\xJ�xJ�x
���̽�/S�8�I��I��I��I��I��?��?����)�)y�ɜ��L���S2�[���H�$<z
���?��?��?�²���),{krRK	ߞ�g��S�²���),{Jvy
ߞ·���)|{
��­�p�)y�),{J�yJ�y.�G�=%�<�eoM�+kI��S���=�eOa�SX��=�[O��S��S���<�<��d^ċ%�5���p�)|
����䙧0�)�{
˞�qޚ̩��0�)�{
�¼�0�)�{
�¼�p�)�z
��¨�䣷&s �&<z
g��q��q��q��g�¨���
��­�d��p�)�z
��¨���)<z
��£���)<z
��£�����_	�ޚ�Y<LX��l|2�a²���),{k2�5a�[�㊯m���O��S��S8����>��O��[���'JV{J.{J.{
/��˧��ZO���������>��oM>O�O2�[�cp���O��Sx�^>��O�jOa�S��������>��O�jO�jO��S���>��O��S��S��S���L�N?��O��Sr�[��W<���
����)L~k2>Y��ߚ�O|W��S��Sx�v?%#>%#>%#>%#>%#>%#�5�x�����dɧ��&���?��O��S���>��Oa�[�ߕ����)�}k2WRw
����0�)�}k<���)��)L~J�|
���9��9ߚ�Y<V������dӧp�)�
�ߚ�Ej�+�)�
�����&s%�)��)�)� )� )� �ɘ�;��O��S��SzZ����J�@J/@
�����&���^���;�5���������&�:VzZ��Im+=)�)�)��)=yş�? %w�59�x�����9(�7(�#(��/�#(�#(�#(�#(�#(��/��/�7(�#(�#hM�B�-�#(�(��/�(��/�#(��/�(�(�(�(�(�hM��Z�����?���/a�K�ƿ��oMΗ>Y����%<I�	�_�������%<	�_��&sJ+��K��v�5�<�UI�	���,��%�I>	�_���p����$���?�597��(a�K��K��Kx�����/��/a�K��K���d��7׫%�%�%�%�%� %� �����H@�!�(��/��/�-(�-(�-(�-(��/�-(��/�7(�#(�#�!&Y�%�%�%����w)�$y��q�!����������&��������xn��_��_�[P�[P�[P�[P��_�[P�[P�[К�E�&�-(��/�7(�-(�-(��/��/�-(�-hM�!&��%����牿H�AI&~IBIBI&~kr\��7(ɿoM�Oj�A(��/��/�-(�-h�+��������\��������\������������������������ނ�ނ����������������d���UҫPҫP)5��/������4�&co�������������������d^��R|MzJ��K�J�J�JzZ�1��I�Bkr��$;�$;��������������ϡ$w����5�x��>��>TI&�%�%��%��%}%}U⻒�ߚ�E�X�+Jz)Jz)Jr�Kz)J��K�+J�+Jr�Kz)Jz)J��Kz)Z����@|R�К̽xg�w��J�:Jz3Jz3J�PүQүQүQүњ̕���k�&�&���?�J�Sz3J�Pқњ��{�%=%�(��(��(��hM��������w��\��\���� %9�%��%�����I�'��%Y�%}%}%}%}}y�,��������,�������%��_�_Q��_�7Q�7Q��_�KQ��_��_�sQ�sQ��_��ߚ�Y�Ez3Jz3J�0J�0J�0J�0Jz)J�&Jz$Jz$Jz$J��[�s�:Lz$JzJzJzJzJzZ�9o���8>�(�(�(�(���%5�����H��H��C��C��C�&�+�&=%�%Y�%=%����I-%�
%�
��q�������ҿP��ߚW|MzJr�KzZ���_IOCIOCIOCI�Bk2��o&=%��%��%�%}%=����Q�J2�K�Z��Rֈ��P��P����"�����P��P��P��P��ߚ��,����7I�CI�CI�CI�CI�BI�BI_B/d��C�oP�[К̕x�� �������&cߐ���^��^�����������^�����P��ߚ��K�g�$w�$w�����?���$c�$c��g��?���5�E����ې������/��Kx�N���/a�K������/��K������/ɿ/ɿ/��K8��$þ�e/ɰ/��K������k_­�dݗ��%Y�%Y�%Y�%�%|{	�^�W_¼��՗0�%�{	�^²���%<zIF|IF|	�^­�p�%�z	�^�%_²���%<z	�^���%��%�y	g^�%_�&c�����%Ly	S^�dΗp�%Ly	S^�9_�dΗ��%�x	?^�fǐy�:G��.��/��K��.�$#���+�#w	�]�l�0�%9�%wkr\�!Y��]�vOa����Oa�[�1�d�Oa��0�S��),����)|�>{
�ݚ��˔��)��SX�),����),�|�/SX�),�{
�=�Ş�bOa���ح���CS�ۧ0�S�����i
�=%�}
�ݚ�>4�ٞ��>%o}
�=��nM�#�Дl�),��5�?�Uk2z��/�gO�eo����Z�X��n�s%9�S��)\xk2f�5aŧp��X��$#�59.���d���$_~J���|�)y�S��)��~|�:�§p�S��)��s��	>���qOḧp�S����\�M᳧��S�ڧ0�Sr٧0�S�)�uk2��`oM�E<GX�)���\��8�!!<����)�����)���z
c=C�@�)<�vzJV��z�[S8�)�tk�yR�H���l�)��&z�\��IOᤧpҭ���f���>%�}J���zJ���z
cݚC�Jj�~oM�J�᳧��OɍoM�C<'�4�Ϟ�?��nM�J<L��[��I��.|J��.|��W���CX�)\�f{
�=�Ϟ�bOa����SX�),�{JF�>{
�=�Ş�bOa���حɘ���Ϟ�/?��nM�ǽ�)��vz
;=S�I��)��\�7	'ݚ́x��Oᩧ��S8�)���y
�<���5O�t��:O�y��?O៧0̭q,�+O�[�c�|\���o�Ϳ�w��y�x'����7��]���O��/�w?���K����~�r��h����ë~�r��/���O��O���g���ǟD�Q�����<�G[�ϼ�{��_>?8�����I���������2������Oܿ��g�%�����}��G�n�?�����I�ױ6'�}:��=���������D|~K�W�~&�n�����8�^S����g��_�\���C���P�����k3�;�����������si�v&�������yh�9�{x��{yi��K>��{j����$����nm^G��Ҹ��fq�Ă���k�%�����Ĭ>7���o���ru����G����sō!���� ��N.�k����?M2/�LK<�m������?_�f�C�_�o��u�Ig��pH�[�}nR�6�?�8���]�hw���@�I���?�Qvi�Ù��Q}m�F�潣��%Ǹv��r�؏�&�7����y�@�@��g�}�~�[�+���=��w|�h|��U���x!|Q_�����6�޼��Q����솲o|�i��|G�'�_���:�N���y��O���_^�o�cX�y�����r�y~L��:�����P6o=���u�`��/Y��A�>���^�)-(��!���绚���������������&�������'�9�W�	�\2�g4>q(߂�7���{���C����{���+����]!W�.��#�g�C�Lȯ���]��z�xť�����s!�`��i9�\������g�O��&�ו��~h���;���?}�h��k0Y���J߹X��*����\2K��/���:d�ѵ��b<���c�W���d5���}��`R	��_]�zd�1V}^)��4�E����ǖ�L����d�}��pH��u�K����+��]�L߷��
E
�Ȓ���}Ez�(低J��ן!�P��Ȣi��g]�F�(��bmOH5J�t�n1����#�Iů[�s�V3�!uȾr�>e�Mq'��;�嗼������1�|����duK������+�wX����7K�k����<z/ꇬLY�!˫�b���~E�}~^��-��*�E.ف|�Te}d��x���yW����=�18ɽ��/���S��\�:�x�5���}9��d�HDH	7�_�)�yd���MVk�V�e��=��n�b��}�Ӎ�Y��s�V\!�Hn����@>)��i����Q\��ٷ=q�e��g�.�gs�;
�6��*d���Z�����(U��]�Z$������y�ҵ����f���ۋ7���嗼��1�.���~�m�e��J��;x+￧����&|}�di�z��eo�c,��Ց����ՄԴ��<ε]�_��7��OɁ>-������#��}c�D�{�vK�?jw�)�3����߶E���?���4��W*�;���:�k���hV]}J������hZ�<e{�ܹ�m���K{YE�����~�8�6�����Nr��xF}��7?z�	�C���hV�(��y������.˖��K�wSU�X.�/��k�8���߰����ƙb�qe��Ly�9��7l�SJ��[�(�AՖm�>e���r��R��/�'�	Y�]�l}ߔ�_��˕�s���W���=�S��`q������c�#�)O��&%�����)Ny�s��Q�c�'G��CW���+�jH�f%5�S�6Gny`��Z��~��o��״�xB��"e�y�i�y�ֳ�m,�~��ѻ4������ﻶ���ܹ�'S�����[�0���8��wßd+�V��<����$�b�������󦿏3�C�-�k�K��vo�!���S!ٳ�g񂍵d����%Ki}����EJ�}K��	N�K���~���p=q�Ͼ���쑊�}�.;'%g�����r`�fN<V�Y�?[���;�rm���sł�_�<�	���Ɋ�]���ߧ��lG�_���%�:�!�U0��;ze)e���m?3/U�+ږ��b�:X3|"e�$�
��s��\��<��3��G�E��{ ��)��[�s���K��������3Ȫg)�{�+�+�*�^|#�����Sb�K��Ia�ؚ��zB�.sB��ړ���H忥$��}.mْ�SS�ɒ��F*�L�:y��ϐ3*�\۽y��:�*�c��2u�X��{�l�}�*�<n�[�1����%�OȒm�<ܽI���'��-[s���Ȯf,#E���-N�_z���ꐪ��GcN�ֶܹ�2���-O1�'D�O����ge�1��Pp�O���5q�+^���4 X�mu�+Lii��6x[8<�&ʓ�����0��gI,�,�}{c��C�pk%�������K�ڲ�y��,`��3��EC`��+��՚�Pއ����^3�s�5�Sl��[�#�{^��n���I��\K��N{dТ]�FL{jE�yV�y����aq�)��m鲣{B~K)��d#�ӿO{�*$���n�[n�/�-��F��r�e���X{�����L`ʖB>Ӡe!��'t��6e���u��:ڽe������Re����f^�)���؆���S�^���,�}�R�֖��'��#Ji�t?Ŵ����e��T�>	�=�#�z}#�ɐ'��\����ߴ&�;�逳�C�3yqu'&�ru�g�veY��f/��	�Q
Տa-��=��.W�iz�eّ�r�ú��g��R��m\�棷�-����L��G�u��"k]!4>�:�����hM��nZ�1f�:���u�|�l�͞�2m�qQ�B�i�}iM<�f���PIv�uH����XH~!)�2�~�8�����ɒҞ���±\��W��K�B��8!Uz]�I��Ӿ�:2�!�ҕ��)�&�޳�,��m><[�&bK]��,W���K?� ��ʃ{�@K�ǽ�T�%7�m�����=�g��[�"��;lNacJ��G��3����;VH��m)���tּ00��'M�ud���FK.�|�>.��ƶ&Ja�ڗp�#�{��p�?����)�����*(ǔbo��}$� �����X!��>BS�tm�>�{v6eϪoжF��s�x�d�}~�r���W�>��z�[��y��_�������k�������w{�6��&u�����E�%�PJ����FV(gK�㞲�S�G��y��U��C"8�Jծ#��Z�T��W�NH	��̈%-�����9��/c�ZO�]��
��3��)^���Q��s�3�#��o��,p$�K�����}�\0�U������Q�O�Bo~��C�S�g�IFq��z6�h�.��vʭ<eC�)��GXJ�RMm��X�0�G��um7F6؟���-���'8By����Ɛ	Ȑ���-��R��l%��؍�ȖW>� �! J_���n�j�ik�
gY�D��q�P���~�f�!뎮��n�BpGkuE�ެ;�Ϗ�[l�2���M{ٷ��i�Ua�ϡ��W,7Ә��ǔ5׶݃+���d����v�w�޻�#�|MU��ik�>��0���H���=*7���$����i=�'���B�=)1��0���t�,�����S6�1d�-�O��R�O�Įŵ��]��F֐e���'�`1���lѶ�in3�m>i��/΂�J+�����l�ȳ�W��"�B�����]�.ǋjJऀg�Uk�h�8���<@A={��z�,�އt�#��%m�v�]�?�Gn���,�L��h�����ŝ,���i�[gG}�b�1NY��O��.��>�4ɎU��y_���%E�N۟�GZ���Y�޼�>*������)�l͕҄�73��+�&ޕ��X�W�ۄeS��K(��/o#�Iȹ/��$ڢ�4��ޱ�a0$����9!��9� ��$�f��'�[�2!%�y�l<�P�mCxȣ��!ǖ��e�ǽ�c���ay�Gb��ro�O�E���d������t[�B,�=+�%�'R��% ߔ}���Y�{��#v��<�-� �5����L��ш<���6@�d��K#�#�V|E��loM����_�-���B�}�#�l{��Z�ҵ����~�<�R����%�Ւ�-�s��&�I��l�Oi���ץ�%�Xeh'�UA�}S� e���V|�x-��S�7��%��|�G A"���{KZイ0�r�z�\BG۽xHv_LyT��M���ʯ��ǐ���}Z�kZl��=�I�}�r	����~u��Y/F�����=+?��b)��)�l/,�m��7�N�9a����r�I�l��$%��IӒ`��6e��4hL�C��������J�C�����k���RH�%�=��[�  n�~]H_��P%+hY,�@����s���R�MɅ���-O����:���H�C�^�һ���.I@�����5]|�=���7=OL��_���9�{F�.�y6�����d���'���g/�bI۟�D��KW�E6��T�,na5��n�R�*Â��~!�����!5XL�����5���X��<��O�]F6j�^
9)���O�[�6��Kx�%q��	<g�����a/�e/�<R_Mj�����ȿ�k4Ũߟ�<����)�����V{Ķ4�K�#�-�@�
EX��y	�����v!�/��}�h��ĳw-c���z�d]��d:MIQ{�r"m�F�<��o�lx3��̑����ҷMK�lK=K����Yxi�[���,nٖ|a!�25�J�����'[k���RD����"�aM��mH�j�H��!!��`��)��a]�����-mk�K���K`�dI}����E�*�+M^���ц�����z� ���D/B){ԂP��5G0��@�Ms�: yƷ$F��W`���C��!p>�_&�$a/8x�%~E)Jm��I.�򱎕io�{�1�C�/�j����H��v��Ӗ�M\r3���({Ԃ�a,�i�q�ͱ��nY=s��w��p,��U��Nֿ�.RȾ`ė�4����
�ҔM��'�gM�z3�)�!��oa%Vy�!�pȱ$�i�4��a�2y��{��;(%��-��@�%5mH+�x$���Οw�o,KV���罹�osK��Y��(�aW�Rr蓻-�K�"���2���=���%o+ _��^6$�2K�S��D�Ϲ�Z�s�~4�����'h���F��^���_#�CZJ�=qx��P �a��]J�c�vu��H� �A��E}ik_�|�i�;I���DM�Κ��Iy+3ۑ��(��K�o��Ų���?����Q�<q�kS����\��	����]Vs�U�:R�e)L{�>���
�BO��Ƃ���Ζfɷz5hD�K����)%x�MǕ=�m^Q~2�/�+��v�C �������tɦ�S�d�}�k�2�@�gN�7�	���#���bN�e	�&vq�^ܗ��)�X����1b��)�,�\_W!/�����S���7����lB"�,!��/hk���n���!��x��Q �7K��gۄ��R@�ۄD�ɽ�Z�ޕ��L��}�'�Mk�����z��TE/��rB��j�kA%]fK��qV��!�����ؒi�GR�����H����Hb�}�G��F��6��^*d�+J�+�o��=�5nM����n���Vj�gh���Hkv����I��H!��Fy=�YK��B���N�J� Ʌ �֣�S�1���Y�*)��<��[�5��=���,n]l���$�~�J�}'�9�ˬ�uiu�(��Ҙ�e���k�߄B�(����ټ؆A�����9%4H'��x;���Vν�A�1C:���/[ȳ����.N��[��F�������C�!�M�ϵ��$Fy��j���\�}���ʞ�xs�8!�T=���KַD��Ps���HK�?_x@���m��?Iu�����s�lҤЅ�< *i��Ѥ�]�^�}�6kq�ҳ$A,�.l�c��7�R�8$���2��vN�a�Ǣ>�%���SNs�cY��,�S=�R�O	/�GZ��x��<���x�e��4��M'��A���\���S{��#������G�1�<�_�#��v��f���5�����g�%��{�$՞�N�����a��7��"����}��[d�!���p��cQu��}ߺ%�kC�:�-fsɲz���!qB�uIl����C�N�K��1$��}b+�di�~��x��"J�ҹ���C����}�����<x#9�M�lh�;з��}*$3\V�#{A�9#{���W��U$��7bV�H'}m����<H��W�4饈d`.���֕��4[[+��5}�w.ٴ���.ݥ(���ٻz�(O�R^}�?E	hQ�}$	祸���}�%�ѽ��W`\YZ�iy�K�S�-/�>��<��H�h.���u&�i�2Т�d�����d{Ɨ�{�+���/Œ��^����D��Ŕz^����b�$��lgZW���x��<����E����.q�e�l^�.��~�m�+غN�(0)�^�I���E(O����菵���-jq���G@�^�>������OG�þ�eY�JC�{?���aݸo�?�������������o������??������?�����?������������������O��?�����_��������?}F���r�/�\W������?η�Ǟ�, 